PK   df�X�xb _  ^�     cirkitFile.json�]ݏ�6�Wʫe��"��z�yh @�!�D5�:��,'��ߏ�?%��x�ٜ�ks8�?g�C�K���fQn��d��j�I��%���\\��͒��f�n�7�Ӈ�����=���~|�n̦]Ŵ�\�Y�ʔ�B�:������:���,yx7V�Q"JV��.*�rÊtY�Uj5�3Nʒ�ʳ���-e]ٖ2*uʗ�N�r��Ri����KY.X�~�2Hj��� ��0RS+5�:�U�1��`�-0-SL�7d9���U׸���q˓ EG��0]G!�p��Y	y��<A�� QO3d}$t)���)4��eV�Z�����뚤��<͖ܮ�̲�s�o1MKL�9�i$�n�<�m�j����MMOD�!h>"Z���C�*pS�4oN�j3\��RU�TP��JU��@���tR-@��i:���)�ZH�*]�Z�3�J�K�ש�"�)�����j9�NA-��X�b/�Z2ש��*��T�2�,%cU������k:�OAM�,fX�!�
j5�A?�4n�C�8t�Ǵ���x��A�+!���i:�q��4�8P-`�a�M�� -��~��C���!:D�!D����M���D���Rp#S�:UZ��!e�j��Nj9lNZF4lMZ�_P�!c�2
&�hlMOE�@�#"�!=D
��p	�D��(h]"Z�z���X�ܮ��X/yU��gt�c��a����+y�u�w\
��L �����p�Qz�Gᢢp�Q��#xMI
G�8�%~K��a��8҈8l�@���0�b�4��&�i�8Z��A1=����c�t(�uU�4qPL㠘v(��*��A�L��Úi;z�2�A�g(ӛ�8dz���"��\��3�\n.l�I.�v���L+�qF��b?.7w&�1�cS��`�t蕅��İ9�7��c�O^iRe�Æ�R����LA���}�ƽ��mh4zz�����B���k��۠��i����K�A��= ��#h������[7�K�T��Cp�i�Ac�nt�\n����-[e��4b8=I��_��+�]�r��h6*�1��)�Ȩ��E�£pQ��(\�(\T.:�"�7zI��8�%q L� �ā0��a�$�i�H:8�i�8(�qPL㠘�A1��bz����M��rx.7����pT�%θ�\�����e����\��\�Eo�޶��Q�l� ��}���ܜ'pT���,��rx.7���s�#��9G��\n.$pT���N �����	�Q���(�����F��\���י�����)�XU&�̒ϫ��O�4�b�Yl��4�û�ϸ�_����
p*9�
<*�h:f7�k�Tgh��mL�9�G�4M0ٓ�5$Խg�hh@�,jLӘ��
� ʫ�4�:�ǭl�2�1-N���X1ט0�;�e��0�)�\aZ�X	<<� �c�cZ,h�ED�lwK�=�qo0��T	�#�O�yc>n?Y˼�TcF�;+����߻�Q v� X�}R�1�;	�#f���#&xw/֫�K�v."���1&ExW/���K�u<�`�<�n^ �7ac�9%x��ɤ /��@z*7���;,x�~^ ��� �ń�×�d�����yTES�W�sV������s��~Ua���' ap��F'�S�2yS�{�A��g�1 %�w9��B����d�(��`��˦t�0�@� R�E)�`qڥ$�`�I���XMJ�H�������C�8����<��ڀS��0��[
�$e��g+�vp�r ��eL���NR�ԟX���dL����}b Lu���+���=��Q�8 ��G=x��,}��5���5xj�_@�s���8��]p�3l6���0���aX'D��83z���YLthD:��:�==�,&7�c���,zp&��]`��S��*�[=`�yÄ�O�����jX�ְ��Z�&�s�!��,��YU.�h��\��|�Ǥ:5�ԍ�`n%�����-7nT;}�i�N�u
���v��-�n̺y���x��ՠ�u5��A]�j�1�}�mEȖ���9�&6*'d�T� +�ΎY�č�o�?�lcZ������{�:6���K㿢�E�/}G�.=�E׎���I-�=L�{֐�|��5��a��My��wxPo�A&����u9����B�7y%���P/PB��3�[Hp|��2�]ߕC��jﻩ�#��}[��\B�o��R�����"ԋKpi��Çz�.�ߏ�^%�KF�X筻��.�f���k�Ŵs���c�豈�E�X��"~,�~�8	�H��_��E�/��"��S���gr��ir�4�{MN�&~�ɩ���79���'������zW��e�Q!���Ӱ\��.�P�׋ec�j�-w��.֫]{p��%g��~,Z�5~�~z�l�LӮ��F�G7nw�v��X����ψTs������[~������em�J�jZP�����)r�2F(�L�n,���f�]� �%�ͮ-6�(2K���r)B&����c�jʵ9v�g�\�(����qA��(�A�S�����g�z�OZ��u��� $P@OL��⊄�~b~�[�<WU�,��zN�d���%��� =�{�����(�s����ė�\b�D/�lw��uq�f��_�Q1���ȳ��8�ْ�ovRi֛�s�t�8� �G��L�Չ�}�?V��v_��g'V�9�K��"vh��:�Ōs5g��L���d��zi���Vi�3���ӬĂ��j^�(D7\L�'o%����(�SAvqw'�`��-��-(c�a���	���;�[��|�~�E&��=�ά��Y}tlL�ް��T��ԔFXՓe�*�JU%�Ҩ%c;(�	�BS"b�>��ޔ�%,��ȠޥH�k��"կ��K���"1RKp�کl�k������F�v,�ڱh�kǢ�����=��ǧ���C��ܵ�j�Eæ�辻�Y�X�M�����߬얞ؿv������L�b�3�pg��V��rmο5�?�Uc,<�fo��Xl�uQ���4S�_�]���ݎ������M�wulG�R�W��*ުɣVV�M���LZ᠇����F3��bsUҬ�y�Je���*k �LԠ�:1 �_�T�5<�,��a��vaB�7�|��ٍ,�
��Rp>J�:��ّ8�L�����v�I)�q*�r�Vq*z�Y�����Ԏj��橮Hf�4%�E���*�<�������n#W݇
��:~��/)a*�����S�����&�Υ��/:�C�ySV�Y�Ǻ���e*e^��^�E\r.��I�*������h��!3N��Q1��Gc�j�Y*�i����5B5"�Ո\#T0��[���)D�*O�9�s���:��9�ͭ�"J��� ]�Țд&�eZ��Y�W�,�6��ZM�@Wp���ٜ9"dg�w_z������� ��!��j�,�vò���3~s\Pb��T��l�V�$)cv�����@֦vZ�n�b.4���ϫ���X���|0����hk
dT�.����_}�.�(?��s`�Mc����V���36\,��c�=�1yx<���1�=Z%Z4���u�=���cf6�$+�{ǫ)>��)���SD񞶫M��h?t̾<>>&.�k�����������t�Z\y���#��QY���3UE9���,P����|�x�C��ޢ�� �$.2��S�AdS��S�|tʻ8��L9��[ �Z�]�q�h�}Kiawl�d¨�S~x�fL]@#N9��h�9g����"��}*����Q�0�%:�B��2��Ј�bq����^��o2TT�Rq��oX��w��}W`��2�0*�^��r`B"h�a���9�G6���!ޝ��^&�d�^�e:�T"%ʮ'F��#{���{�rT��x��c�GF�O�,��΍���S��9��8 �T���UH�t�1�������QQ�s��^ YB�P���}�B ��Eg� :�M `�6@�dq8~���;Ļ>ÉR�ә?���GÈ��`0�q+��Z�hBjʽm=*�`�4�@l����;�C��d��9��pv::���L��2*�`\����8Gp��3RT@���g��q̲�0��
3X vo'6���;�������a#{��sw�@3���*�4�u�Ug`���0���P���;��4%8���."��[<�6�uTE��	�2�+ ��:(��t@�!5Ԃ�][�پ#�p�h�"��
2#���wMH�l��Y�)���#Oy�dc��x8�we	H?���#Ny�r�m��S�ç,ݝS�O��L�^^����w����F���$%Գ��i���;<�;D���g9<Cd�/sݷ`T�$�02<�qdT������{dd�ϯ����=_��� Q�������B�]yDd��W�C"#��!�g:{��p=dxddHU�bb[R�Sb[���{��ز��|��бe�������"
�M��@ڄ�e�Z��.ZӬ��.yp��u_V�5���f_��~|ݚ�;���wO��ߦl4��Y=oZ$_�PK   �b�X�H2�    /   images/17766975-adcb-4bce-a273-4a591672b910.png��PNG

   IHDR   d   d   p�T   	pHYs  ��  ��F��   tEXtSoftware www.inkscape.org��<  �IDATx��]	tTU���{���JB��H����(���Ӷs�>��n������\����e���rfZg����E�dI �'��m��VD�@UI}��V�{�����WUWd��+l�zsWaV�A�&���Ա�6K�
��9͆�k����qmE�M�th&:�d����d|Q=+E�i��Y�ڈh�ɘ7�����ja���:�|kq�C�)ƫ�'�m�aӅ�)ߋ��:o#��yI�!EA9�j�#��q[�l������
��"	a2n]�?�^�n���B�%�t�*��+������������x��y�=�)ܟ�PxP��e�.�1]��C�,��
���}�TG�/'r=7r���`ܷ������K��*��y�n�IWJ��͚�S��+>��ȪK�h�I�����]�?\�a��!��',�o"|Kѱ�tԻ������VN���K�����ɭ�Q���b��Ah
z`�y���/����#H���)���(pI��ֈt4R���w ��9�ĄL�����T����{!G�?NY�B���F�:�� <N�j���z���?�Zy��Ɓ�t$�&��#�m@�'��5蹝Ɉv����F���^�mm"����-}ʉfiw[�<:u��Y<�o2��s��z�$���~z�g��[M��Asȃ�wL�?m��cs���ikA� iFi���<��!�ɸ(� ~?�s�&mW�Y���o����K���Ha��� ��������Ćj;�\� ��L��e�n鷧z����?��*�����W͍_$ᶄ�u��zY����N�T�\��L_�O/+؟����N��:Rɠ�p.Z)M*짛y�N��ˬ��yKq��݈ʖH&^��3(�Zb��he)�y�/��T����e����������R�Ť9cf�������%ס����fp߃SZ��i�4nxz�
���i�y�k�"���乼`?HFmK6�>O�e���6��d�Ҍ���F�8�(GV��*��7��t!��C �����9)�vJ7�*�HO�a�����rf��b,� �|��Q����ｺh/��4�
6.�9�����6�rW�#fi�����2�?v���/(.��!�UH/W���R�O�e�d:�_\>�'�����Lu~��^a�N}a9bZ6f��?dbK�AM=�{d�pPDJ�sg�w_ɘ 4#Щ��zx�C��U�F�!������
э���8���_�NZ�ϐ��ᛂ�9B�m�m~Y�TU���v6��>�Pu\�޼�6� �}�PU���t.�����ၞ�PR}��T����ܺpס��R�K�:��	WΤ�����@u��LM�Ec�cG�!l�W�#?�{d���r���`�ۺ���.�-�Ң�N(�yE-�<i���;�N�a��)ퟆ�ݔN�r�T8n�T�%�%{���HK��/�Ŝ!��v?U�%踓��gJ���i ��8?�k�IB�h�ӹ��[��2d�T&�4�L�4�!�2����N}9M��Dx"�5�Q���x��:b'��r5��&>߱̦��:��eCȥ2�h�}Y���:L�e�0b��,� �fN�5dӿ�
�%ſ,�X�l��4�J֑��Œ6���[+7ȶ��7vL�f$?��!�֮�*>�Yykȡ/�?\&R�)1}���[�leۂ4��A�iË[Γv�����i�i����?��h�J�t<6Q�����`��?p�e��4G��f�&_��4�41D�w��Ji~�c��=ұ�p~2n[	ˊ8]��j`Y6��t�if��߯=DQs!*[S�W�]��ǵĿ[;�7�`�VB�Z&��T�i���(s7N3L��3��~ |t�'g���Zu����hx�+s�_����@
�)ܕ���t<��|RY�,��*XJ���J<r�&Mn(�^��k��<E^�#�fҦ�.����.ʫ�c��͔Q��+���DD�2aٰ�(�z�ue �%�R���`�Q��l�ƨ�s�_ˇ���l���(KO�����o������8Ni�G/����$��3�C8��6"��x��B��nhC���)c$UD�ᰦ�+*�gm����Z��O�Ɗv�df��\��@u}�F�����1*[�$�@M��������6��$�0n�d�Q9�4Z�J����z���BT�~ؿ�.��Z�8,����%d�F����
���dȼi%���i�Hc����ý;�]���<v���5��_!;����j��)��0淌I�^���;�G�Bv��d��fz	j�ڰ���� ��KŊm�1�h0���G�����������L�cR�r��_����ٟ�1� ��'�����P���l��MuL3��٩TY%2*1o�JKF�WÁ�Fh�χˆe����_�A9����H�%m��s�L�f�n�H��d0��
6�^C���|���Mxh���k��}t���QMu�t�F���6T��O��b�v�aG��3�Ѐ�u͘l:�RY���E�ihF��fLQ��� t|��uM()� +��Ɂ�rQ\�G���:9vUC�?�MP� ��6e�u����ADZ#T4P���*��&�����q����p8Ι/�x4.��Ҧ\<|ކ�Ӳk^�(ʖ闣����
ß%�`��L]�K죇�^�^����^�R�$P�A����MA��G��IY�:��_ʵ��+,�/�B��J��u�p `�`�}ƊU.t��&9\~g��JAsY&��z+Wq[ZZ�眂�;�il�e�M���;�Φ>�_3z���-��Cٻ���A-I�|u~/v�"�����tMA@�����&�˷����q-���w`��J��p�6���6�k�a�d��<%l���`&�s ��SH�U��V�{n<�{������DHNv����}�eH�A�&"�������^�D�F����ț��ɉ+J�:��F8��:�߉�]�R�B��	���F��e��c�smM%�9����%��3���5����!��5��9�w�	BB"�\��=�>C���:��ν��i��P�TV�b}��-Ӵ�ZK�!}!�S�0�=�s����w����m�9B����8I�.:��$!�%	Bb�!��g	a��";��(�iB�QK�4!�xӒ>OHXK�'���0�)���ē��B����O3�5.^�����~C#V��!�%L
?ĊU�+B��XV�~ұ��O��P(6?���aD}I,~��_��08���o	�D�?�m�ؓ�~KC�"���5yz�ׄ�7p�t�҇��5!�h+��%� Q�*	B"`-���*&��3x&%<�|���-��>�J�x<���93]	B��sm��t����s��� �0�H9��+A�	������N;�5�x�1�� �.]w`�f��CA�?�؉���4�q���	�e���������Gu"�ȑ#���E�F������$w"$���?k�W ��#%)/�k�(�J$��5��?B�ǃ�Ay�m�v���B�	z?C����~����x������cw�o+&�X�0�^�����k����I&X��|�?w��֫��b�!.'(*�6�A��!5o��zz�:�+\8+�=�C�mIƍ�����>$Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $� ���n�Qb8i���tu"�\�f�g�y�B�Pyw�.61�e����28����jD��sd��I8�^$��M�y#_�>�7Eh��׼s%oYj�����P�WR8\	������Z,A"#���ҳp:�lGE��T�� ���d˲<L2���y3IEqe�̅�>�,�媼�0n����7�O�y�B�m)�p�0�Y:UrG��l_�k�C&�m�j���x�o�,$O��n��4�N���M�q��m����T�U�M���o������^���^~wa�
2��xf�r\S��'�JR�Ť1��ee�͙�Y�ÛF�Lyp�|��g��^�mQ�@�y��k�ދX��?B�U������� �17���]����p��v�s2TM�"P���|��y__�>�^�%Bخy��W�}���[���[�]d��7t���������>���K��[jw{�h�Y�
ϐQ1O�Q���v���l��d����>D�Ͽ�o�?!B�:�!My�4c�5���٧Y~��*�N�ϸw��L�0����fd>�w��T%2tem�~U��틧f�*�q���>J��HM��c<�^72������h'�W�+贻��~Q��[������nSx_\A�֒RRM�-"������}ءq�![<:=��������"�8v���Ɉf�x�8.��8/����~1�������"�"&d�b�ff�����;F
iŧ��?g����*��Ɛ�^~�#P���{`0wp4��KՈ�HF��QI
��;)-��Ϭ���
]u�$�r9�\(LJ&��6zY1$��H=usű�r:(�p�֦b*�B������Cض�c'�8�e�2%TP��ߝ����Ք���t��L=��2��\!?�xj��#6�T���'�вa)ڶ�Z�'�m�ʗȎ/J�8;��o�x�T�Z���'u��l���T�mJ���'�I�����q��a��ߨ�G;�)��%�'�PB0�08g*1���O�=���ɮ�.�"Ye���Xv]iIt򓟙�0��>|��Kh�"����Ua�3�Y6��.��B	�-��1�ӪB��O�dI�v��G������$�o��:���2a�<4y� �ڷخ�� �HJ�p���ROv���,Ƀ����aZv�Ŷ�����Sr���N�<��Gvn����ww����#,�$�c�5f�	���}#����	�Tג�񹨕�.>��1M����K['�^x(f^\>/n=N��$9�<:��NI�»1����CXOo:���pݬ3�h�IN�c��|k�
~��<w�2*X�z~N͒�%~n��"Ҟc_Ǣ|%_S�_�q��|@0����g�h��&m�/���;Ғ5�*:��U�)AG����x��9���82;��^L��Q�X�nc^�b�����݅�2�*,3Y�����n��4b�
wf]�����)d�&K�3A�g��l�����XP\�qa^�ՙ^?;|�8������d����h�},���ɸs��thn�k��̺�<ɉ��|,�f��l��_��K�D��x�    IEND�B`�PK   6d�X�@M��  2�  /   images/1a44c3f5-ff5c-43a5-9e5f-4b6f5eea1ee8.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   8f�X\��䓝 Wt /   images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.png�	4�k?��)�RB�SȔ�M��(B��"2g��ls�Hl�D�L;��"2�����d�f��:u�����}k}��ֱN�y�羯�w���~��sAI~�=�0�ֳgdT1��Y�N���O���j�~�;u�����*�{��-;���gͻ���w��jګY����cp8�uKs;�+���V���d�=�~�Y��#F�ͭ۩n��J�5ǆ]��_*^-	�w�s���b�_����v���O�oԽjV�kw&X�]g���_}��z�X�C��Cї�J��EBxU~?X�<q��8�][�����[Zvۿ��C:P�}`_���)�V�,i�)G몁�{k1Зs�-�9oo����׌�i'؅c���u�_���rO�������9�n�ž�#������HbgO��l4��7���N�/R�
�PSHJ�M�+j�g=Q}�O0���+�j��nvl� ���4�3E�w��|`K*�t/f�ש�P��n��p]C+{�QY`:o�|�'|�݉��	z�g�����vL�ݮ2�	�$��86ױ7�x���-mk��\���9��晭��`�~^Uj<K�7�?�Rw�8!��f����s�v��U��E]��,�Ε�m��O��]�7���:b��c)x<�L�Ѝ^083ٔW���;v�<]<RUL��8#\����IY��+o7����촷�!Nf�O�Ń���2U�7Y�9����?�O祣��R]�G�ǎX�6�\�O������BA:/U���1?�z��^D��ޛ���������\�A�:X�����e�}y2����}ǩ;�n���:ś���|��j
��.T5�Xv�@~y!l���z5��8.� �� cdC�q��m����F�3��F|p��(�tm�~� ?�(����A0>�^�<C��Q:�R��j�P�iN7W�����9}�n��8w,[ ��s�Uˎ����b'c�����l������s�8�>e����<�=��\Y��N������/���ԥ��j�ɚ����V5�螟�qF:&��t=;�3�%>_ �S�Ҝ��!;�6Mn��%3�;�=D+/ک��d�G��Ar2��v7��gځ��n�J����O혳h���4��&�ڲ�i��^�gj��z-��G��Kh����RH���ak硲9��
z9wM�Aj'��A��v"o�_�-�
1�m�}�����<Š���!$H��X��^���1�ZJ��T�I�m;��x6�~�c�5�����)QI:k?XS��RK�#��	Zu�0չjY�u�!*�Bn0v,\�1�5^����	)K2
Cx<�-�p�c��ˉ�	�4*Y1��E�e=���;U��`�h(��+c�f7�LI�{qB�ez_%l�²��"k��ǋ$̦Bٻ8��pt�P���M�#��Y�"w��1xYYr���� Hs��\Z���X�< Lu\pY� ,F�$�����Ǻ���<*���(�ZMUAY�hZ^��vB״�*lާ�����Mv�]��* w4�I��*�H�RG[�L�:��Y�QmY�J�s���gy��e���A3= @� �ϑ�#I���� 6�����S2)�i�8�ɧ챓��������y�^$���v#1u�vf�3w��(٢�l��,Y{�I�G�~���+���_��&5e��H���p `��k�k���E��v���H�V �~9`���Saq�?�q�l�2�总�>K�Aj��j�֭����d��M��u� �:2�:)��q/��H��	 	l *��?^���uލ�ݽ�:r�,�W�w�t$o��^�ޖւ��B.�#����<�V��zd��Mr!���M�H���wl�5�p��3:�k��-���W��M���룔-T*u�AfA#[ǳuz*��G6pw� "��j.�R��L�$6z�XyFuܱ�pg'w���:6�x��̾M=�����c[�7�r�\��S�,rW�Q1�A���K'Ɍ�\�l)�v٧ᵜ	(��s_p4��$�/iC��X��ZH�^m�{�QCt	�Oի���NS <�eb���ʸB�V�!Z�8!sp�6&<4$��BH_A_br4��������I��i�
�;���8��͈�ğ%ƾA�J
[�z�j$�7B��7�_�"Mf��nkӭ����ddd��4���ݝ���L9ONM�lٲE|��R�=<<,�R[�1���o�+,���������m~����\�v��CV���Q���"���6�<"�����!NΞ�G<�Ǐ�jL1��ٚ=��������E[��������������1 Y����+ Gz�E�<��;PE�)��ƙ��H�5��=z�С��b?�'vk��>>0���]�>`/��k��X�?I'S��]Ix/�_����h�꣌bL��e$�\�x��@�k$�q�s���v>�4!'^���n���F��@US���Eg�p�W�fA����go6�H�J� �9jq�4��fWm�� �k,aNԶ!�e������y�`���Z�$�%ͼ19���bt��3Uԡ1hРq@����Ψ�)�d�  ^���Al�Ν;k-3�8o>V�hN?H.�'gQ
�Eqs.��i��Ғ�p�jG�X��N�g���8U��\#	���KJz����9��;�#���@�E�TiY����U^�i8
y>�i�$/�����0���� I�PyzUM��	<��Fm�E���e��i;�S��cRl�bσ�Q�������8���6�|2*���ZQ�n�`�0l�����	,I��=y�M��3._�R�Ԍ=�g�^t9PXI������*�IYj�>��Ǖ�;M�;vݢ�Χ��<����`bbR]"�4�����c�)����)�ec���/�w<�%I���ݽ�dJq>�#��ґ�<�F���b���}'҉\�F�i|8Ŕ0!�C>�ȮZ��X������V������f(Ɏ��i�p\���ܭ��X���3�$g�BlF��D�.�jm;������H	�)
�W��DŇ��T�V�W�!	�F {7��t��6��f�8�-,�FHyH�6�\A$9�TL�u�ac� ����Di;=��Z!R�rc4 �G:v�\#jg�e�㎝	��6�<<.&������D�$y���#�/�)1�Z��f��J�$9o��t��h ��ǌ�sFFF��s�k3�\�@ �� #�$��jdO�#""LQ�=� ��b�g��ʹH2���>�TU�ep�J�� QwY�8�U���g����˙�R3���?�"3����X,Բ-�DH����	QQ�a+�-D�����A����qN����Xl8�k�'��E�9Ոv���3�m�D/�� ,xq���a�
�ny;�}Fss�L�ԒQ�4+������P�	܍��ϴv��b���}�I�xgr�%1+�R����nSBb�e	S��W�m�989Du�C�V�aB*v����[)�}<6�-Ķ݉�cccg>�0(**f��4��I���,͉�O� t�vѳ��J*X�J)���ik��>Y/�1HbZ��o)�*5u�j%Z)5C�����ȃr��z~)�S	�B���[A� P��2[=�h~܏������F�̍ёX��5#ښޫ5
��w�n0#F�|� ́��{�T��d`�eU� ~>��L��P�b�gڙ�kn_^���7ؔ���X~�Ƈ�\���T��-sVf��!W�:(ks>����q�d����¨ց�6[�fT�$17�j��W�;?=�+p�����g�n03���J4@�G�����v��� q>D������h}=:���,��;D���U��d �L��m�=F�ə�/�>����~x��3磹���[�NQڲ'�Y�&kIa�a1���*1��k�T���Q����6��=�,;J�E�N=~ <r��s�{|8#g� f�����!@R*�ut��/{��|�ȶS���g�<9�$#3��\���;5wy��K��~�B��Bv��x�N�����.O��&k��SV�zJ3[�u�j�=���Z]�,�ϫX�^a��<�:����v�I��Q=�Qu2_�b ���g�v��ܩF�\�fPɫ��F����'��ë����gff(�ε�E�l�"�`;�5�����&ȁ�� ��[�	t�9a�繓l�S^6XX8��X�W.miI7.ϴjϙ*�='~4����+ęS:F4��ɿ�ʽ0�㢢����;�O_$���I�ւGORKlrE�1����W���<˰WĲ�P{�rJVX絅S'�tA��	$d�ѐ�dAJ��8��I#I]�#n �n-�	�����$YC�L�\�~����e�8�u�#��ܟs�z����yd�'$�R���bm9k��*�E�.�i'���Ea[=�Y�
Q*��\�m����X��rFm�ER�:ݨ}J�
��B\����N������]J0�dF@^Z��<�ӵc��__�~Q����X�B�`cx�2�^<��	d!i���PNM����sʀ��^�l�)�.
K����x�%B9�i���@���D�Dzm\R�O���ag�e�>@CߩOCM�M�g����)����3y��m������G�{����s����0�4����h�
���G$%�
��T����ܜ���O:����Ú
ܒ���N�/
'���r��V����1��C1O�+� ��&v=	�{'M޺eKխ�:;��F'1ya�-[���&����ß��'�K�:q�s/]f�D�X��S�v�s~�\vr�|;%p�B�­7� ���m�O,���"�s�ԛ7o	�������+���4d�ڨ555fm�9�c��J�G��֯_�M��E�:^�vtϾ}����A��`7#�TF@Q��S����y���=�ss챗��o>�Nz�$�C'Ӳ����0�Ķ��-����m�z7._��@v)�#9�<kЪA<�B�Q �s">˅H&��L��e/q�؞�R�����p��T���$� 9����u�@�d��(2�5/Bsꌱ�:{�����4G'��ƹ�)]���)5{6n2œ8��"�m9Cj>�Jgj3��DvT�Z<��	n�'�l�[X�ȑ#ۣ���#]�o7�޻�O�c���(�S�|WWן ����ҖM��J�UEؐ����tۥ��l����0?������nU��r���A��,����F�\�u���Q?<��-q��ݻw?�j˪@Y��;���:sۓ��C��$��V�'���}O�h)����Y]���qJ~6o�����=)�Ao��,7�z3���2 A���[�:��Z�p��H�TEIy$��;U:�0	����d&n3��ff����
Od{&�2���98��`3s�J��K�y��U�.�H��͈�1���v�5:�����`�T�չ����mqP�ggԌ̖m� ׉o0�5Nr��gzק�����i<^;)��q�-l_�"��fc�8�N��M���)Ԑ�����gTK���(U�	n�aq��ԟ)U��.�����`������4�Q���aWb��+�J-x|ُJ:d��*`��kwp򕗗��m����Ec��<�iJ'���Q���'�Gӝ�l�+¢�I�V��Y�(��0��-W�g�fc_����Mg9�@����1���E�������i��6 .�����tcE����W!:���(��B�D@������k�=�w����#P�rM8yU�3.�|(b�YX*	u�)X��qC���>̯�s,G��FI�:��Dȉ��Q�ns:�=�:Y�l�O^�ڎ�����^���jh�w��A++�P�kj.�#nB��y;S^���d�"��D�x�GJ�I:Y��IU�>��`v\تc�ÇUB���)�=�����ŋ݀u���,P�(�d�$���\�/���1K��l-E �q� � ��l/�R�q�"���!��Z�>.�NP�v�j�����T�������SM mGZ�<P��8���S���l���M������FID8:5��p�2.Xlx��*�a��M��O��
�V�[� ���PԱ1�c��p �$��q&��q��&��h!���=���3�>dP������P#ܔ�0���Es��S���y' �I�\���.)�c224d��`-		G�}��Ճ"m7�a>\�f�cg	�bb-i�^|R�_-W$��3���Z:�ej�CV���Q1\��o4Wt�E��v��@��%��?�4�T��ͪN��-$$�cU]X(����I�� �������;�߁�Ѫ/{����og�E�=	�{z*�"y�`Uh�G<�66��mV [�9o\�b�>|x����aaZ��Qb��h�����@�F�+q3�E���lA���l����,�*�DG�bo��h���nŽ����J@U�>r�B�w����,�M=������7ɘ͡211]��]����Χ�%�Ǩ�L}����'j�|�II L����(���[��C������{{��zP��)��v����ph]��t?������e�� 	//o�ҁ� !�|����q�N&�?y�j �4�9��9h��a51솢�¤3�ŠY[�m�]?|�g�柵׊B�tr��X�U����h*��`��3�{q^P��R�k���Z�z�p�l��y���Z��r��pe�3,�����NV��)UT@C{�W	�R)cmED�O���Y=7撮�ˠ�A��K��j��e޽��6n�7h����	#�'��4Fv,i�4zm��&�j-�n�˩�,�Ï�B��\��ʌ����?{�������N@�px�ʝ1!�>}���=_������=�Ү��۶�'�����)���p�\'��I�P�	k��8�:5���E�ha!o�_F��{ �P����g�Z!�=E����l������\
�]�KӁ��������oߞ"���x����LLm)!�ϐ����}dT.t�c���:�� Z���M�n�v-~@�銥%?99�4O�����~ļ���(��)̈S����N{���hǉ8���� \T���/N�^��y�_�����nC��N�[�1��JК��J�� �w6_?�O�LF�?PO.����'��V��8%F��9>�1�Ɋ�B�pc�<(Z�rnٺ���ֽ��I�J^𖃠*#����C�ub�j/�������e�(����G%$X��yp��L�����f�Cx�8<��ӓG,�M��y��e/Ī�ܿĿ�dm{K��7@M�ww����p2{'y>���#���=d���Y j>�\��'���Ă�K��Ǐ�It�MT�i� �>�A`�i��[.��;� ��$���X8l�d#��SVUAPT�����iYY� 0-5�r�BuB� x8�j�n �QX$C���K o ٴ��+*+��f�Z��`I�����׎��?`����W��MR��+�~l̚�趶��!3���Y�] ;�N��ʼb$?��Ag�����Г��l��?�z�T_�F}�Oi��'�'�Ų�Qg��� F�}$���4;�d�SP���" �����Sw@z(F�O�<[�!qMH2@]�����0��ʣ�K�x8p��h�3��k�,}�rT*A��Y���w�\�_or����xb�J�B�� ��J?���k���Y����lL-Xt��FTpD�&׀tz�& ��'UQ�qh;�	h�JJ�@,YP<���s�ű��e�rvs��,Ǚ��T�����)x������}������������=���rg����3����G�3����;��D
b�U��	 ]!=�JH��7�������X3D� ��~8s7�cqH��J��!��`���a?�-$(#S���Ufk��F��ƭ-�S9']���i@\
@��I���9�)�f� ��-�B�)�.�� +�h'�|�ce��.�4�Z�=o��u)�!Z=�����kI��tx`Gyz�f�$�9�q��O��烍w����'<�"g��(t�~��bB`�K�Z!�f�eW+�6�,1f�H��c����l�\@�*�>���R�Н
$���T��J<�}�:�>M��##SV��a2�#�Y/%c�M���JW)6�b�t����=�^-���%D�"�»<@�j��}F!6]\�4�P�d�5�l@bdd�3�7�O<�r�HPsIU���"35��l><ߣǎ]���3+�Ft����H`%ϣ����Դ��[�c��r�m���PPa��S.���v��%t$]�#��[�faf0jm4.����x�A��̌����cj>WE��)@Z�]�b�r��1�j	�.z����+Ϡ#Ц4#�a�۵[�5s�ym���7+��V3�<PdT�;6�0���NP6�F�2�,���� g8ņښ�?��"2�r�ږjd�s��ʊr �#�� q�\#�\;����� �+�k5�h�`�f��B�'i�v+7L�]��P}gn�H����}�e�xG:����i����?f��`N���X�^sy@AP��d���*����0(�>1�A阮Q�د[��.��q���TP��H�gE*�A��@h�ĽF��{��2�'6T���]sV��*��~��H�0����NZ�;������U����2M����ΫW� ���p��.E�i5B+ְ]%4��T_i'�!�b��]7 (0���\>� �󮬟i�W��qi=g�E�^�q�F���( �!h�Y���$�\��O#E�*�̰>R�[74�@����r�Yf+|�~��E�C �֤��yތk�xߜa�*rګW�XxWO���?��Z�m���2�z!�;�ǀ��qD�$Q�%W�p��F5c\Y?��[�d�������YQwKWk��������Ⱥ�$w	���Yf�LV���gavR�m;�[>��"�'�ycw[���� =D�[x
Wn�ViH��y�Z�<��h^Y���/;4���V�R��E��I� @�>d�~9`坹�t^v�����::@����l�㡆�=Nx�{�V���r�Y��/5����-2j{�7h��=���x<����ͥ/� �,��m���	�M�����W�3�o]+�S�����m�Ė�I�I&�ϙ�m�D<�y�5�����(IO�����@ 'u
��r�	�+x����A8Y7{�P���~�=��+�3�B~ et#xǩ;T��qǔ���e�MPCt�|1p��"0��HS�ф�z�[U~���D̢�_���.?�l@*7���|��[1䩄�h��88QQ[�n���y�|*�c��XYEq��nP�	�|��w���9x�1Q
���H}�Q	���k��/--� 'N](x3�x'@>��UTTMN�C�"..�{��fl9��*ׇC#��vniYm��l��8y��zfz�)߇?�2��;A9�I����Lgq֞�E����-�/)u�BCC��9o���I�z��n�Kݞ�_�|�|
�?�7$�]�Az̺.]YX�X�<_'6�F�L ����<~q�B8���Ig�,�-`$ɨ�ŉ��iQJqq����@�؎��)Gq�����Ԗ���t^��րw��8�7Q��6��>MY��W�d$�[�8䦵[66��>w�ꞯ_�3�Zn�[~�߉����ǝ�:*L��?p���-��O�s����d�ۈl^�	�ݔF��	)�1��q7�*T�LdR\�B�wg����ygɊ�>HډH]�v��q�����N)@��b>�VM��y��F�q-��@͌|����UϠ&C���G1�����w�7�w�7�w�7�w�7�w�7�w�7�w�7�w�7�mÏ���+���_��/o葆�ʵ�o~F��|�ESV�V:o�XsH�=�t���B9�=�����6lHz�v�'�D����{~���)����=�v��RG��e��î�:{�]��f-�0��%;�����e��3%|�*��6K������"֦�A���A�+����f�g���҂mn����*)�`3|QPSW7�aq���B۲��͛�ʒ�k��y�-��L��v-jc0Vִ��Z���)uCA�	S�^��%�kfff���i���/߸r�GP@�bu]��]m�F̘��,	���-..�222.u*���,Y���^rñ����@���?._��[�YXl�{'���;�ܪa����*����H�pC���k������u�p��`���-~�V�,�I,v�oWHn�pȀ+4�"]����� �q}A���ۅ���i=��I����c��sh<�A�:�\����+k����=� �Hc��?Jv�����*����yt��n��
���ޖ�?lC	-�Ǯ	����v!(x؋��θ��(��R���:��NP��'~��!�`-&��L�$h��ӋU�;X�쾵���3g�A(��8va�)����N�/�@�O�%j ���2�޽�Qq�QK��1E���1���)��驩�SH�s}��2E��񟹛�j0S$H�x�Cg�V�����#R��d�z��d���L;�M����ۺ`���跉m�R9<�e��^�-ߡ�:i�4�?��4W��|5�A*�˸��K�?���rER��ݱ~c�*QUJ8S���ERػ�}��U���ޖ�G�M瘯�|�ʍ��y2��y�E��LV���#�����:u��I��ډ�i�s����EDJy���Y�QuC!�g�Wֽx=:�\�*�i��0I_�#	����V���o���5>_�81��p��4�!?�S��c9X��u�٦�������ee���l�2a��gN�="�i�Y�mF��ڪlV�b��}C|�;�9�A����J����zV�/A�/LM���&$�i.`�����]d}��%�k_tH� S�o�ݧ6�����eF�U��0�t��t�Mf�uq����l}rfh
v
.\w06C�~by����D����v!��.���ɭ���t��o�i��N�<r�R�d�6$"E?�ABfTf��ej��͸%H������KVD���<�)g@��lw֞�C��_������fi�0c��4s�)x1g�;��o|�O���ĝDov����F��]�Ѓ��>��Q`ő�lwמ�EWT����g�Z�����u��'{��y	���U�]=�؉�I��=�Hi�*=�I`�
4��]�=!��Hr���.Խ�5��5;����#-��� ����.��|K��\�dD�[�Ǝ��U���pڢ��0~n!]|9������}��D� bM$�]�G���=�=�^3�ۉ%��+�'sǻ-O��-6��߉�{8�b�h�9M��]���EȈ��D����ח���WO�hz_��-@�?�>5 �/���-7ڞ�R��A%����y��o�7�	��3��7[�}��^?|�e���H� �|��Yki'��E�_q�,��>L��Vi��AL��0k���y��h��?���|����0�Bj���Ō�Y����k�:�Өb���t�+6���aRR��h�G\��%���"=���;����ͪ?��޼yiO�݊��Ҋ�-��E�g6���f��C������փ�c�!z�d��5���bXc������׈Ý��	��M�F��d��gZ�)� �D����Gz���5��]w�A_���e�����b|�!$�n��Gi���U������Ⱦʚ|���n\�`?5�m�Y?�f-}��ҫ\S����]�(���[¿4�����ٴ�8�0!ˏ����CBC�/�V���-�@��_��Q��';��d��^N���$c�IM����AC/������Z�n����h�
�`�v}�|��zV�0�1Ӌ��O2�"X�/�o�j})X�=E�
�R�4Z�v �ێ t���[���������@�^xL����6�з!r=�� ��I���`?"��R~�،�@��yet��� 3WA��X��7��4���8�yZ!G��W'N{�ox��ߒ�#4
���l*.M瘪���E9�0�y�S{/,l�K�PU��>q�g7b�B뿒�K���Z,Ɠ�o�CƢ�v8����"�%^;��\HA���NV��8�E���U8�$la�^EP������Ѿa%$g����F�K��&4<��3���{I�`�����x�e{�
^>�-PN��nf� �E�����f������Bl�kKِ���Y�i03P���@+w�-ETr;�����C����"�}Z\(�'�S�*���|=�8���8��1�S0O-`#hm�C�h���2�=����<d�B ?@��˒��!Q����ьO����_��N"�3�xF��N@����]�8#J�!Ǽ��a��&u�M���&�a�,�ؽ���8����+���g�x(��� Z;��m_��ɰ�E�s���T�>�u��F��.�����z~ ��L��3#d7��������/XA$��?�lTc$s\t�B��뇂�
�����l@���މ��h6�l�H���,e_� �Hl���A�z�*.!�|<<<��
X�q�3�0<��^�%qY�u>�Ve�~ڪ$�Wۉ���z�w���-�MuD���pɏv`Yu;��x	E8k��)���?��N��X���'��m�-�ۉ0�4gUq<���	r�����3Uq��F1���� c ��X� ���ԵkSa �����;;����ݳ�0k��Sؾc�´c����V���D�����xy�N^�Ի�EZ��;㌔%O)�	��N7Y���oO�U����\G���߈Y��%�	�v�*lEl�?�GE><وa�H�����W��~R��R�3��B�z���$7����
�������9$$1�9CO��J9��k]� �~v{�b�4��f~�{x]��T�(�f�&z�����Ca��h�S����Ok�7F�Q���>'�a��������WT�e���2r;�b!08މ�æ�p�̨h�����V�x�O�ڦD�Q���׉��e--O �!E�B��h-72Q��w��/�Ϯ=�� �sV�y� �e��ˌ����ՙ�ӛzC)AW���I��Y�O�L������Y��.'���3}�YP�?�Z�ztz�-�S�ML6��h�_�n�c���c
�(��iw��%)����?�*6]�t�h2wЎ�f@�����=Ok=�@��9�ݿ�?��X0���I�'@?2����Մ�b2\�l���'���O�O*4Ґ̚���j 8�z����;C:�5\�+S^E;`� c�����#���]��=�v��5|�#�(���m(W�@x�0�R��1��5�݃/�Ճ,�֞�p��$>�as�#���7�%�a�n��^���/#	'M�ȯ�t�C;����͠
V���^ج��E����<���b�6L!݊�~�˵2W�����6H��gP�@&�M9-^T��F}�
]�	.@Nd��}Z��%��܄���Z��ap�@��)C!���1�q��YSQ��*��[��?�mï�����5'��(A�i�VYPq����0�xƷ]i��WǺ'�#���E%���S5u�G؊��k ��l꿭�_�����?�%t��Ŀ�s�Z��a����������I�r�e�X+x F��z?-���}���wԕ�cl�p/6����,�	�!��8�l;Q'�h��Qv�j���Uh����2��<�M���v&��	�;s ߒQO��X��j#7���]��U����0��wOm�4=�����`i���Y֟ T}�F�/����&�� b"�8Ү�7��X'����?�;*�0F����$����b�M����^���i�$u?@�+hs
���M���0䈍Ϗ?�	3F�[�rG}�����f�<o�iVmb�����THV�Wc�9��I�+�@�MB��&*r�aRqd��3�{�H���^$0r^~�p V*7k� 	�or\ʄ��O���?es{�6���e~������Ʒ��G��Nn��뿭�=N���n�\���?�٤4e�9�\c^p�4��y�8Ū��%c����Kg��ˋ��-��;�����Bl�O�+��E�?�(�O����7�����@�|����\���`���t�k�"��B�pƟ��iB�b`������b���wi�ؒ�=���ڵt�dt�=a�b,m�ձ���6� }��t�Q- �������~���y�ٲ�t�X�
�w����ٳU�� Ԍx�ڞ�Ϧ21�����_����+`S}��*���0y����ʀ�̝�B�1T�C�H+�<(�ߝ宸9z~jd��:\�tB��c3�"���#��9&HaY��:�,37�ߺ���;v��=	�;��J�F��Q�H��V
�8�@{NA�G�J��"U�]eF��� �?^��Y�� ���E�>����˔Y�B���������6=qP� ��]6e�Ώ���T}d�݅Q�/S9�IIg���i޻W�[��0�yi��^[�سe�����e�d 8���b��>��%�nZȁ:�6  1�v�,}"��s=�hž��J5rNt��Kq� ��\!��?����� dd�I�O�ā#�ոVW�݌��6}{Ȑ�$�e��&C�d��kDm�Rȝ���ϊ�
�������QUvU��j���9�
T�;f��Z.���nnn��6櫒[䴑@��^�Ƹ �4pgn�
�*�J`>ӟ�Js�2���8 �)��1��ᰧ�"ȶ��R9��d+�@m���&�����	
\hLq/�ٓ���������jO��P?u�T�SHE���0���g�LH��[�n��sQ��ޮ�l�u֪`(��gn [�Vо�Bp����DdJ4t�1�煫�2��L�3��pUm{��.2��H�2�X��M���c�<�'1����Z�'cPu8=0���ь�Ʒw�w��L�����	D0W���!�&��ڙ$u�V�+���N  U��z8�[�tm�H��H����'�ƨ%�x5��؄���w��F�B��X�m'�B(&>^��*���P���7����J����������m'��[?���^�D(��t@z_mq*B-�YW��,`����5f�@Z�G
SFRؐ@/!8�ʭ{���Gn�WK[��fڛ,$$w �菲1�cD�����������5U�^�O��3�/D������UоO��P����iW-��	��g-`��d�;�NgR;91��,D�7��@hѤR	��(_�籽ծ�����՝+�౐����[:��#<9���0��=��G|�?p<���A0���v�}e�����|�h�D\=�8�E:tv��i;��7��'s6dp�;��1M@݌a�c���\�y���L$ᔦ@c�3mV9q�1vA�M�I��X �"b�WD$#�oli���vҎ�
�R<�n����#t�	wa���C��g��cUrW=�����ݨQ��Z#��*�h��?��J`���Z�|k0��bW�L�'0M��o�<���/;��|�k��&N�E��e�_}��ĸe���\th���d�<B�R�2�!h#��85�� �!�WH��r�W�ov�`��=�Z^�A���hU��� >L�>ubK�x�/(��+��?�X=#C���~��������=�ʓ�r������{1����>�s�yT��DtЭ��r�>^;����q/�^ϔ�q��ؚ}��3��[SY�8������N
�0���:�!�3�ƽ���}��Wδ��c�a��,����=�&݄�ak�f�w� >����-��Tsɂg�j-�l|k�J�@�Cb����ɓ��❄Jx���w�}�o�s�؆�[K�33����I��T��!VV�Í)P'?=��U�h���!#��� `�i4,"��E:�ɓ��6'Ǟ���L�b�?��ŋ�����[oͳ�GO����cos	$ݲZ�B��|�.`X�������ۂ%�9O)�~������6��8G���$�V���5�T�����G���B?|8KO���=�m������������0����`́����I�:�t���-�^Γ\��'�A>GOh��x�����Bp������_s����Ir�&��;����߅��{�<���[J�u&u����@V��f�̈O�)++��8��K[�n��ӭ���q��^�V�B�!���ʁe�8hL�����S{��{������H�����2��NDXx��z�|����s����>���5��/V~���!�l�~����S��+]k�?�w%�+�	��(}��gbbb)(�P���6�����EG]]}n)+F>�lr��>��%��Y+�@x�Λ.h�a-Ɠ���,�Nd�d�-���]�1�|GD�f�>~��#���rc�A�ׯ�y���!���NNZ�K�����{�u��rT�>~T�f��2Y��(yU%Al�;9�Jo��v�1#����37AY�r7�Ÿ��8���A�+w��r���" ۜ䆸9BE�ǹ:?&��9�!NNcu��4j�B��wM
h�N��ᚐ��-���c��~�ߟ+d���z'|���'���=o��);�[@?�^l�A��n�<��S�R���n��Md��Sԗg�{2�浓q*GCoGw-+))�O?Qu��ө���ߪ�㪳�����a\������!��t�ik�3Ǜ7����(rssy���B����(�JJer�տTs񨬪z�Գ�q�����Ruz�p������e��_0Hi4vw�gdd�z��IF&&c77�	�A�������_AZ�-,�~2�iΰ��:�#�ֈ$���x��~�x��T�^���hj2���P*��(`�)g����%��� ��?0 vt�PXD���C�)Gu�8�c�i0�Y�vi�7�n�A^[m(���?����DDD��3L���:?d�VCJ��t���cg���V�E
弲r9������\J���@_כ���g:�m�w�^��k1��e?մMdh_.��aqqq���f���#�CC�O�ͽ�8a'WE�r�)�\���
Vr(13��R=e�F��d�G�,��a��O|S�kOP2�Z�V�<�Nk�K[5�\v�Ƕ�ՃuJiP̦[�s3�t��L-BnEۉ�~��U��+�\LoF�T��@���/hFJ����x��������#Y%��A&~�{���KcC���Ѧ&;yUu�;�gf�NQ�O�g�n��M�.����F%TTW��d�k1��`�-����'<����ɹ��E��1��_r�q�Q+w�[.��E݌R!����=����$2�ZU�T 
a�∦3��2	�6��O�32:)�v��M2T^��Z�q��~���=�u�i�����`v3�c䲚2;��^�0���C��S��]O���
iY?R܉]9R�>H���8�A���S��E����/M*��<e�U��jZ��ϻ���S���{{+���Z:�����t}ӌ�`�L��i�z�ܦMOOW-�9�r��o�����LM��l�n��3
n���B�Y}���gز�c$g5٦m�w�>k%�H#E���>
}t�!ź��lfƣv`0/~��$��ݖ�b�E�:�Dzgj����z2Z���<`ဖ�~�ݓj���@�C��~>����C;(Ox>���<��R�A��������5��c����W�l�>_�I4g�G�3���{ߌ����CQr�E��B����V)��ۂy��p�H@扐t���H�N2���d��d�I�*:h�i��_�й�%;�a-<+&d���O����o
�ٚ�\�:Q)��B��I���޶l;�Ź���O.&4T�i��c��W.]w'��#�E����>(��\x�2�P+��.�	[(�Ap �������-o���P��ȳi;�t4������om��n��k��c9y0%����G%-����\�
Ni]<��A]���e[�� ֩%Q>��:t)��u�o�	ռ��(��
ְ�����Ns�ܝ/Y�Em{�y�*ɺ��@Q�wE��X�s>/�Ͽ#k�D��r�hc�ƶ��i���\OV:�ݧ��2C��]�2��i���i����a�|~~~^���N��Zv�����!����8��y�����;kY�k�jѿ�P��ᱥtH8M�aX��w��$��!A�б�7�����+`�/ �S�'Ӳ}SG��������_��w���N6 �W� ��Z-�^k�AҸN5h|���3���bf&+�:��8Q�q��TT��]䧪	S�b��J����5��i����=*"�	��7H����%%����A��c}����>+fRqɎ�1ݞ5��/5�e���`C�*R z3lv�{$�Fm�O]y��)��)s
��{�����'�u��W�p���rK2$^/�
.�i�+Sާ﷐��2�Ӗ�ҝ��$�w^,��D��^����W�2�0�k�H% ��?5�R��,'�t��,4��p�޿M������{ )�]��BY�d�*�@BH<(�9��f6̤*H�|j�Ce�Y��(�Nj�Q���{���a՞x}1%���hK%�^y�u/��@��H�ר�h~՜+�uJe��,��v����	NB֜p����3�(��7fW9����zí
�cq�ҹ����䅅힝�	�	�|��1���E��SEZ��)�̳c��Dvy�����.ԫFF1�[b�l�v�sS�G�X���5��W}�	a�VK?9�hU��$��@���@Su`,�4����M~�x|�k�@_��IƉh�u�O@�$9wƲ#�[MM��/m!�	��Y���7�҇�dd3���qcע-�8��7�����΍��Uy$��wz(w�@�VB�x��ͪ�g�����fy?ub�t� ��s�ý��S�aE��+h�w�\nll�KH)x`�q�%�P���#�.GiJt8
�Qr_�6%G�3Qh�V�#���$	9�PIr��1C�c��`0��{T[�����w���Ƕ����~�����z�.(u�|ك��)�/�NW	 k��6J��c������w=A�p�cgQ�U.���ݦ{_�;M��^-��](w}v@S.�"j�M%��� �`��Z��e���ʣb��9R���7�����������p�F	���LM݀��]�v1p�l'��2��( ���A�«��6	#�X��|����s@�+�33o���6zs�-�}_nn��'�ꩾJwU����u�ӣ�O�6�9qh�t_���(��<hmG+��d��M��8 �����6����W��$́���A��3�L��~`�+n#Ң��M7��@z�5�e��$�C�������kc9;[=_/�*�j�<(��lS@��|�v��A�я )$0Z�P���]��`�+))��5��n����� U����-?6�*5K�%����h�Wy�T�N|�� ������^rT�U�#T����Jo����_��Mml��&h͕�X�o'�X-�\����/_*�G3?3Q��SHD�F������s]�
��P=&�S�f�r�=�Z�_�1���վ�S�U��!��ʀ�9 N��C{�*�X|��2��p稽�x��ɳN>�\Nb܆������s!�W57���>
b[��yKPHzbH��+������=7��|��5`X1 >F���MuP@�.���0nM��ﺲ0)�24�_jȝ>EQ��wt�{0���±��Փk3�Ï�65�ݱ2�$i�'�F�������f�ʙQa&��� �~�^���q��O��?�H���R�P,W����|4/'⩒�(�j ��=o��-�9��K�@�W�
L���dq+��E�� Xt�$RH�<@��Kq�Æ<3��&����8�י��ك�"IӼ��}�+E@��=3����f��/'� �a;����S�����c�`i?���w3`��w����Ɩ���A(��P��
��p���>?�ذu��##e��������r@�
����C�W,�%�x��l�~X�oɅ�)�ߞ{p��U�#���"�� �e�,����<ܫ�>�M��i�'�r�q ����K�wJ���k�������4��jK=�>��m�)��o����jeB�G|,�����i���������LDc��
�z���H��*�l`��V�Kh���t�m�&�[�����j���a����r�\ ��QSS3�ճrF�^�~;�Wd��C�7>P�[�6Ƅ7��c�<����=��O?�pKꮟfHi�� F�{����3쵑�7�����
���Lܟ�|�;��U���&�������֮!��ݳ�.�B��%����^By+!!Q=�)ǒ:�h��X)�N�gx�yۯF�y3�^�OD��l�׽������ӿu� �?Nr]������G_&���%M��H���W�E�%��W�ߚo�l_F�f��p	)r��<�	�nj�u�'I'癙��/m�z����YJ_����+��l�F�����ࠇK: �U��"+'e"�p$4� ����h�j%���6*}*�kf��;s�V������|������q�������ٶ���{)�Ç���e�t���T���.�~���w� NIx��F��<j�������&����/:;?�v*m�w�fk[�f�����U����j77��t~�� 9��q|P#.��0��e�}����/��������W㱎��D��� ��y���U����:�����~[�0Q�NA�rV���#4����l"��^VF�dd��k��W��VY\,a�Z\�����s���蘘Ѐ� ѥA�(I�jC�հ}Y���{hٍ=.̖�$F'߱���Y�N�Dۣ!�Î�NrO�(������v��YϞUG��3��qp0m�RF�B-����r,i�V�����â���Ϲ> �����팭���0 �����������Ǫ������w����u�u�PKo����Zb����q]������+�n�9D��;s�� "�	 ���k&c�OI0 3�]d�X�q���U��Qᵈ���
~`x! �)��������@�ƾ�X�x@Z@ԓ��I|	�c�I��
9Q2�E~G���g��#^u�]F>�$"��P�l;Xn[+oy��q�V)��"��M�v���N ^��v����\��?�Л�ivdۙVB~^p���LY�l݅7��ͽY�L�@�����^���Bc�7R"8�\��� �^��W,-U�c�ΐ��<-~�ղfN������Q�RȶǲWwӪ���/f��>Tv�(QWW�E�b�W� �󯶯����i��a6k��+�I�f��WW+���-et�U?~�1��c����_��-����q�3O�:����7�����g�эc'����2�xڟ��e} Wn��V,O�[����c����˹�?��8�>��`��� ��b0\[�:-/�;Hs����={��i�=>L\!j�{LLL`s}� ��8{��[CY��|�.�7e[��vv>��Ѐ�G��T��X�}Tϼi/U�5������vM�B���n��IHJ��1uu���z ��8��x`��L�ĥ�=??�{�g���*������� ����u����8G~��[ /�����"��j���%���S���VJ���N��/�yzYK⪪�p>��^3ccO���۫fffՓ��%�;��۫��ҕ�Խ�[Y��o@��q�e	�]�|4����D��/#���6�����Z a�06�{��nLxF��i�������������ΤaC�E��e�nF�;�Ӧ�1zT|��9 ���\7h}|�� ��RލM����7w`jzz�@?�x��$L }O�>%-��"&�Knt]$YBL��u9~��U΋{XYYP��=����&`d��/"��I��	`�?���}�����nf[He��o���F`+Ma+v� ��]px<>Ɉ���K�<B�q`X0��#-��i��뽯|�����e�&l�����d��W#nm��Ow���ǹ����9��PW�(T[������֓��6�Ү��'mO�ʁ�- {hc�+��ve=}��*T`����{5lb�����^+ݓ�[Tص�R+�\�4��s)���h$�3��V�(U*�����E^ɫ%!'c��e je�;4���C�+�h��w�mV���>cu��D[�qkMg:�K���j�������g���_�4����8w�!N�oh�144�n�[��+s7 xP�V��6�Z�Dx�Т`Э�T�r�i����t�z��w|~��s��iƌ7;y�4�6u�0whge);=ee踻�5թ�8
���ި�+�v��U����a�k���a����i�\���=,?��0^����������vO԰��U�a��b`-�l��*��~������M8j���}�ڭ��%P�ζ>�mQ�& }\	윜����҈���"	;00���6�'V�b\Y�L7�u����$Rg�`ЋY.�_nW��g	zYՉ
>������믬?�_H=z��kȱ?�v�0p�K�12-�r��{\��QT(�`DS�N,l�O�Uz�<�C�'��g`[ȏ���jD����]�=1��E�C��U�ʬ��A�m�J�°�2I[�.Q�5��+���Ñ�? ��P�tiZ�i~��V"�K�֩gX~X*�X`3U��1C'��Wג��5��h3��_ɢ����V������x�����$t��A-֌�a�����:t�q1���2$�4�����A_Ӕ�l7Tϵ�4� �r����T�Z#I�� ��n���-'8QJ�����m�f��y �I<��m����zY�IF�@����~᳿H�L*���-�HG {?��~Z�Ն�
�2�3���)�7��"z��T1ޅ�CC!?mF�R����V()B""����.J���`��{ŁJ�J6^����M�~�n��b�/\�<T,���bfb��άI��.l��jj��l��j�&H]GҧG��1xY.)�+W<��"H������4���f��"��A��?Wn+d-�(fM[�{��.�\�25�f�E��Ti���������8�y,�@�Mx�$f�+ɈjЍ37_����bkR5>��u��m��<�
�";V��}�x���
�*�����@{�0�W�]y�c�ka�����
��bك��e��Z(�H^��;�8��ڍ�{�H�XL_mp����Kֹ���0"L�7��>6`��w|�͋��[+zc��C^����T�?v7��j�7����}�ƨ:�c�j� �܇�&~�#�*=���n������,�����s+�d���C6�u��T��<����߃�9�Z�C����{�>��.v{ &H-��+_��I#-�e����]��؈x���'�n=�<��x�^��сw^�/��b���T��4�.p4�M��ivv�����v�e]��i�&������l޿,8###�H��Hٿ[�� ��vw�y�.N��d�m�l����'"��m�D��ӳ���2A���`�&\MQn��u�����ۍt�ID�`���$���o�Y��~�����@���7.�FE�5=Uɝٰ�9�{e����N�V�4�b4Џ�9=�-�-������C�~�L���Aph�'��@�N��S��aO۟Ys�̙iXu���N�Q9�i������Y�1����x�ǚa咣c��������[��b������8�<f>���?�\¤=��/ޔ�
�����J�����W2�0Ң�:m�ߩ�����K9����?5$�U��>�E%%OK��I-�x�3,��6��mؖ����O� ��2h��T�2"����8�~����c��hn�%_��A�Ic�H2R��po	߳�Y��V֋��xds\��ZΕ�Aع�EM�y;�k ��-pѾ�G��+�����KkFA����xGx�J�c�Q����p�G����]�i�Tv�%�N��ی|�B���=W/��œb�(�߂o�e��wl��b���<�g� \q����S~ʖ[���d���3��cr2��Z�0�}V��YO�֙���O��ˢۄ,ye%��:�__��m/u��-�?��v�"+֒94�+�6Ҁo� [*�n��Z�	@�@�J��ه�R��.���S�!Qu�����������W�7??�1�-.�Yي����nR��9%mR6z����L�)��-�H��+���;"���q+՚~D^(��7߇)en�ҍOP��>����[x5Y�:�'2�.25��.��m��#wX��;�bE��0�5�&�#�*��N�.��.��5:.��;�蘹q�!w�G���7�L*s��>١�2�iԐ,-�4Y�f(���`օ�w�~ȵ��q�3Sv����;<����2K�{�:�Gh�&j�)h�����U�@�D����h{��s8C��Ʉ��&?B�K�dr|���q�ȵ5�������mx��һr#�{�k�;X�@�iv��f�����������]�Ƅ0�jc�:��z���*:�A���@~��ʱ�ӵޭ�홗��t�����f�<�+��щ��%m�G��$bJEn�U���a0ڼYj(V����T�r3���22��&ƲH+퉬s�@/ll��}.+�N�9��&*���&�<���ɂ=��V)_/��tқ��^fH
Zn:�W*B�`����7d�7�٠��;/\�ȐŶ�r~>�>߽�ǆǟ�n���`V!��[E�z��U��h��Htt��
Q�i�a�3��8BtdQQ�0zV5�1@��B��n��f~!��0|g�p[I�R��<�_9� b�BF�7��1�ӗ������c8$�0�E�t����=��mV��X��vޏ�ͲME-����ЧvX;�^D >m}s�m+����#�ye���T]n�Y�y�b�Lk%-Vu\�a�s��^��p.wp�'8��8aQ�K�1Q)��NS�0���O�踐���Q���h{�2�g��#�k��0��xهk���^)U'��ϯ5[*'�����ʣ�<�{��>�هߢ�G���P��g�>�Y��%s$�c)yB���Ǘ�8q}\	 �{"EY�Q]�(��#pw�_���@��6��K�ei��O�6����+X�e�_ȯ�!z�7��UQxݨ��c�7Û�en�<Zx�e�Y�ph(C�����D�N�&�3n�f�րi���o���!ħz�ge�`dԈ*}���'�>�݀�sK�$��m�uy����NΎm��y�>,��Wceee��_�d���\:�ٶ-95u�b�n�	I�+��iӍ��}�\3�;�ofN����l{3�D�Tٰy����ƀ�nG�$�ȓ�`�����o2G��_�y��{�_�ٔ	o����{)_O��L�ԌN4`y����u�/8S>��!�I�i�'���܀��:�VC�*%W9?p�7�gwҡ쒐q�\O�0�/��X¬�^�Y x����Ì�̹+]��������I.7��
�	����+.*��"��~HkqX��,7� �`�n����=Oڬ@����'��D���p��� ����c5���l͢R�V��S�*�Dzκ{�g&�������q=+횻��2A��;f�jO���	^.�+�2Z��}��E��)��G+%7�_v_�A-����{�����i���6l(ߢ&B�T��@�U~v�nZ��		'~���E!���5a6R�w#s@ڇ�]��1ap3�N^Xp���6B������*՞��:::��*��ܹ��[�X��;�^�E� �^����k!&-�|eHA��!h�X��ʫU��)cn�&�`$��퐻rԅ�MI|?Ha���2I��eц3���K����!}�O����0F�	��H+8H�,u�������b�sA}��Y����m�L���8�0��.����>����c�lJ��'�O���	=~���V�Y�|s�Z���;Xμ��9P;� �:^��n��l��͛7�����V�<V*ɩ�!�@rE(r���6�Ti@,=WC+oۣ��=�E,�/�~ɪekWQ �]��[���q6~	HE���tV�_m=9��p����L{��r�^� eq�9ϑ�bCa5��<��,6�lGe�Uj�{�XY�}y���$��=����jӵ��g��2���Η��Ne���f����nΐ%u1}�j죩��(�@�*݊��;��ک�
�(��s�0,���?�}�(�=��D<6Rn�aP���㉚���C�u�z��;�o��H�����M/.&v��i�����e����⟯8��+ 8/gBj��W $��:(F��.��=��:���|�%�T�ϟˋ�����#�CYv��z��)���6O^�
���0G��`���FG� �G*Nͪ��wX8q��V0�ޱ݃�ʈ�|y��Ju�H�G+pMdv�u��H�Si*�2/���2��=�o�^�?bo_��D���n��+��nQ��Ω���\��.=�Ep�C ��dF/4$i�~f�� vrDffT����������i�ϱ>|a�P3ݰF�N����{�Hn�I�7*�p(g��/�����l�n�F�X�oϟ?�02b�I����#Ms�N1}4���w�[8lk�<V���@�-�O��;.��U�����, �;JJJL��^���O[5]G��w�����(����������=�tD�H���nU&ˢS_7�G3�\r"�^��y<ձ���4Y�L)������!w���g��b�C��e�~\�0	�������>-�K��-F_ �+Q/���樫ѽ�F�׌�����A<=zT�h���prМہ=����q�.�F�<^����T���	�39�L[SЪ���^Wn�VSq�V+u�k�?:j�^�q��x׉0=�X̌�ޔ��N�xw4�%�	
�YEq���E�u�[.8%b0�CZv*5�f���R���||,o�*<edQ����ճ�.&\܌6���h�0r+SA��ڊ��V�O�y�}�?<��w~#�����s�*�"��h�=�VQ�X:�����PKK���Z0Z���jx�t�!M㴛8�0�g�koވO���u\4r�fld�>���Z��P.=��ߡ�ߚ�i쩪��
���G�役9���p�I��펜����(���"�圁�9���ۦ>��T�4t>Џ��_!�;T���X�f4=x��`��U������#!�(:�@'��"_�ǣ����|�M��b��JQ7S����5�(�� ��*�E����w'�����G�3�6�"�!>��#��<[�w��;�+J?��M��@�r�S⨧Ib����u闊���P����
�B�Ǣ�bG�� E��iSx[�ا�Ҕ�\�>G���䭘=&�^���+�b֎����
�>����JZRR�*{!!����_��!U�m��(�_��=9���q���� �k�~�^�Fss@T.����k��*��@u��k `��m,첤�X��^�r��+Q]��0��lt˩\,�>�}Db�$�ƛw�o�	� ;���uU���#zyVf���Z�e����	��t��4VzW��gn ��fKhM��t�)s���zXI��D ��P�x&�ު���+��dȢ���Z�S��<�5� �t�=��?���$\����R)7wd�tJ�ˬ�)�;U�mD��1���ۭ�W�룻j/:�[������CIT���Z>�Ϫ,j�c��M�܆P���+��Wn?����Db:K�Yy����Q�&�f�R�N��{�A�ǯ���!o�0�����@|�;���[��d2d�X�d6ڡ��q�����Q�^�&�q���<nP��-�����ĸ�].6�ژ!��˽�+���W.2��p�\&�ٜ���W=qV=�A�y~ }y�(]=i������k� 6�[��'�+��#a,�i��1�*���
�zU��PF����FA¼��4Z>�q��C�z"Cb��7�Q!��.�Zǅo��PUU��;�z�8K�q���9+��l��^psJ]���R�dB�UV���+�PG$��b���|[5�����O4�}v7�oQ��1)����?;SO�27���ӿ!�v�,Q/�u=�຾�I�QPH�)�����Ԭ%�LX~U��ϐ�S�"�o�Uy�F]Y&U�V�#�s�:�����ڬ�ʖ�� �=� ���P�G�z�b��e���?��o�lq�h7O�(�=�Ͱ���R��M�ڕ�d��I����С�Vi����8C�	.�W���SA��A�������G�v�"E�(�/v�+��pm��ۃ��M�J䌌�bcÊKn���Q���lRO&��$s/��L���VA��w���r�ƒ;���4�ϟ/�f�sgwT��8�����8ӌ�<$z(w8�m�]&��m�J��莠���3/7���4�WJ���kp疏8L�Eܳ�L+pd1�rA�.����ͨ�Y��'�7͇d��/KE,ݸ*��Z)d�)��MGG+�h������شo���Y�����1AY�����Ύ�u`�|F�k�!ON7`^�J�Ga��TC
K\�8{&�6"�[HĐ�l�jȦ�i���}0���n�I���+e�R;gg�~��Ѯ&�)༓�qZ����x�AF�D b*w�</�cr����|�L��<w�t��]�8��'i���=�Ya,��z(�r��x�R���:�
�^.&�l�Ϧ��3g�<4�a��^�|��޼�Wc���0�ԉ�)Ms�N����Z �7�[�ܽ��M**
��4&8k�.�L�`�aq\Pǁ逭��o�_9��fl~^�1Da�(�^GUu޲������D۵;������@�uB�'l]�����'�֑���fn��bΈ4��5L���w�Eov���^9YYM���������8~��X�-7rG�w�[��%8�T������A�����6�C���nd�W;�r �W��٬sY��_�KɲV��bHP���ԥ!�n��n&�[���Oϣ��I'�=�\ִ��
ك��.,���K@c�>KNUTT��݊0���´j�V+L7}�r��~L�߯!��1u��Ծ����%������d�v8
ݡr!]�� �:rL|8^ˎj��l%���� T�)dz~�mO�G>���S��ǸQ�&����<��	�#�(����SIR o��;h\����b�}r7C]nKU��a�����t����:n��
B�!�XK�@�͟B��,[q�P��3�v��*���L��X��Du&K��lrH�wG&��#�o��]���t���'�k�F�v|=��b?9�o�0�"�>��k+���**���D��Lfۦ�q��rn4���$��[��/!mmہ�|5��� �\N�B���������f�%Cc)�.O��yXT$e�̌��g�k�%��*���;�El��k���#��A vʄ�����MT���R�j*�VBb˅�vK��)=L�=υ�%s�|&~�lOdsd`/A}?-eU�v�gqH�� ~⢢��D>�������i
8��һ� ����rcGly���!�Թ�[}A�\?U�	"�Q w�����As������6g<�-+�����>;S�lB�6�S�����y(U��;.�m��W���8y*D�qM���X���ť���D�����^������ �O��9|�]�����S-P��ϡ�J:c�)&=x3^4�t�*��oq��Nĉs0��]�O��ݝ UgT#>�O����G�����̚<7K7��Ik�B�4���B�'2X0�j����z����>�4"��'
��^�#"�/����X��b|^��d+P|�ŋݟ�uw�b�6�S}�2��?s�V� ���!�"�}��ޒ����KE�<߀o@��yx�l��k{�5xR�c	Z.6Ѷ�'��鱸����7 S�f�mo0�#zY^`[�%��)h9ڏ���/����ע�K���O��hT��>��B������;�ԗ4W*j,G���?W d��`�H��Cst^-�������S[{5��q��9�+�ֆ>�X�����8��Ư������MLLJEx�.��������f�	Qt��7��b
��j~!(�����`<�tz��"$�d��fD������[����%ee����P�lbM¶�ē��p��gk�[��|		��Ç{K9I ;Ҍ���B�߽�f��R�O����͟?'�8��ݒoz^،|�n�:�I��a�4}�H
Z
>$`fZI�_�,N)�8�f.����֭c�ma�Ʀ�7�GF����ó�I��'�Y恂-Trꮷb�����6�~��,��H���_x<6kh+�kե���o�y�&��8���t�7���?�0���+A��� ���\����@�����(������+d���+����(�OK�[����<_f��� ���W۟�2rJ̗>0�$J�����@o9�Q��;jz����"����D�*�cW�+M���m6�:��Z��R@���������z"��`l�L��Y|�9*Xn/P��gn�G���<ϸbSO䉓'���-�v���ܰ�?ַ~?>g�8𨷶����d�/��� W�jb����������b� �Z�>¶X��f}���;s]��̺�!<�:r͙��~����Z����
�vS���>��	�!��3330cL�%kq̙��6C�������x���Ѱy�zu�x�����I�s1F3yZ��
�ZM-Gю�����fTdbC�5��h93���ϕ�5-7�b�㮌����U��������Ji�dhW�7i���r����ap���&����cR��}X�*z7�>tpy!<s\��ł~�a�I��H���
a���-�cd5��Bjd�cЕ�6�u�۰(J.*9'��v��_mo����FX�s�˖�#�+>k��n�a�P��#�� O/�<ŹHr��:��H�	&	7�� ���g <L��N7n<�3�A����5�S�Q=��3�&9��Ϙ�1g������/ͰK�)��$����y}4��ڼnT�e�A�&�^n��-NC2/vwW�^GG�x#��a�)a���}E�Y�a����O�GZFa�jt5�&����S*N��S�N�v�|� �@�����8���/�������]rGY���:T����]\9��kkR�,���߽��nH�Cr����c��W�C�����n�����:N̹��W�Dϵ�o��]��CNT�.�# +��� *��v���d��&:D2�c �r�6�WgF�
t�
M&=9{P\��(�RS��^<qQMDt���@8��s�q����͏D���2O�ډV��˺�5>:z,�2��^#����	�ߐ��'�x����X�a�w��.��:HnZ�Bm�ݑ���9����#UFC��wz��368��ZZ�v��b���%j����/pU��e���}�2	L����)�c�$����O��O�G(�`a:!|'SW˳u�S��%Nz�r!� �����w�HB��\�x�0�	�(��\A�����W��湐�kQ�˿l��J�x��_m��r҆��l��D���_Q�z�щ=T�!��5�c��&�I�q��7�x�pQ٨�D}*�iҙq%Ǫ�sg����۬$b��8��9��݄Z���u=�J�˗o�'�>\訂���$�;��'L����i�-\�,uö_\��Z�����
q.:�d��i��Dp� ��W�)Zfðm� ����C��_��I�jb|�==����rpL�w^�.|X/K�_|'Y��ȁ�4z��&�m`�ͨ�ɟ�%�
�2*6����qh��<�����E[
�ֱۆ�����v��TnOA��F��Efcf���	�������5�8W���]揦�c�`��R�~���M%�)�I���`9V+^�E�<�����J۞gR��<��g@����t4���5�N�[�������� -���ߟ4���y�A�œo6[Vr9P��.#<��3RX�L�E�7k��`�C��5��I%����t:�G7p��_1��X�P�������9�/���zB t>�~��A#j������ƋO�&�������"�$b���Z�9����Es�u32A;�)� �vªr��'���)��А����+���֗j_�My^=�	M��r�)Nk��
�*���+q ��V.��/�u���wA#)��!�9X&�~qqH�ԑSW��l!���.&P8(B���8��<Gw�_ǁ�
)C�t�k�?�;��7]>X$��:b1��oi0đ�I߄o4���o/Ӱ��!��#d��!-8Q���������)�ev1��~Ր��"J�[V�x��E��4���bOsg�U��뚕8�E�8Ҳ���p���XB�J����ţ��q�?�ú(Z-`��8tnK���&��G���mf_�.ĩ�}��@��m��P����r�L�lkD}�%g�}�C�_�VR%'��^+��7���n[���	�p��;�M��D���g֯�*Ӏ��ߓsz��n��`�<?��éqhP+�{k�A�_�Prf��%�T��|�l����GLu ���D�����ى.�HػYF8��!�h����R=�'�(�A�b�4J�5~vK;����;H�&�|����bcS��<Ǹ��i&�,S<��fxbe|��#����#�p��씦��ێ�1��X������������C�:IAS4�>��O���h��
��N�_��~c�ܤ�e�"�e*d��� y��#�o���U�B)����`�óS$q#����v�x��Ls��h���[86�0133���>���I�y��tHd�3��L<uIޅ���d�ȗ�촣W?l)q�������p��{���1�p8KS��#��V�b��[���t O���!h��Fs%��(
������a�s����EU��� E�ݻg|&��밸�I*�C{©�e��leVK�����K�=ٌ��x4������jW�w�ͅ��&A�J��ٻ��^�cklld��e��uSv����Q���7�^a�w�g`ڵ�H���8�8�S
gz�{e`���.���/A�e�o����h`��sku\���ZT���~YO\NNN
�,Ox��NC��u7r�(����r���9/H� �������wboųQ%�.�ة���
��h���P��#3sK��Q@�}:, 8���۴8;���e!n�S�v6���s3i۷��&M> n�[�D��}��[H��J\_Sa�_�؎\A���=��s���sr&k�}9�P�/���}.���cR��ܑ��"��	V�@��(��l5��5��CW��������V�:�l� )aӭg/�����-W����+0���n1Q[�ES[�9�u��E��������J����dl�u\l��z y�Y�ؽ{���L�E�����?�,a4�̝�#|0|n��6m�H��^|�R��4mȾ�>��V#�~jJ l*w�X��ڣ�y-���]vU�`��)������	*��ʕ+�0��"{Y~>_������7'Ͽn�L�E\l���0>��q�C[6f�5B�@x�_� [�qϿb��{@*jp�cWُ���#�fv~i�#�H ���w�G�*�&T��6�6,��3E�c���6X���ci����-��/Hv��>�s�%3�;]z_�=���E��yß��p��[�}5����K���K�k�`�9�_�aC\
 �t�Vea(^[ ���a�$<֑9�5,29P���7�a��`�훫�a{�U΍VA�F�=�m�|�����K+��?��U�5���V_ m��͛;3Z��� @��ȑx����(z�\�B��t<�%�z�iWp����<���z�|���E�����z�`^�B�V=bg2�C0���KDc5�]b(�cO�%m qy��KE`?[�����}�Fdς77�y[��Bxy+&����X� X�Z384�����oag��IK�Z�lׁC#�g�SkD�b�Kf���d�026��f3p�
Ѝ9%蟕e��7x���W��EM��Z�"L�JlA�\ZUޟV����)�8����j_El=������+0�8#΀�G9aB��'�4Di�PW�#g��{�z��3�~�Jfv��"�ɘ_�d���x7M�`a��>l�$J���6.-�hjj6}�5ð�S�:���)R:
#�u~'w$�dPKK����d���ߖ��*�<������N�������ͩ�m����:NS��OWi~9�j`y�k^Gc�qZ�z��c�B|-��̻9z���kg����s��TCNe����}���;�§zN@~�tY/�ꏀ� )b��8�H�.�<�|�1"���"�}�O��	3��{���/�X��5��Jj��2�ߘ�����y�1��S~l,�����������u���m7y�����S��I��Z5�6^�Gs����'+s��Zr7V��͉;�P�l�T���4�\���'3�i�VqqlWf�M�xbGǆ�@��T��1��o��˿�,f��as9v�_�5.���w2�I?��1� t�N�oэ�?���1�[�X��2��-JT���>:��z������9��˚�菮�?����;��Wް�����a����g�2���\-���.���p\�V�n�$_+誱��X1�����=nT�����E�;��:�އ�~���/HI�,��:��!��M˽�����<�!�<Z��g�\
����<�>��k��-�#f�݇aE2�s�k��L���	;�p�m_�9�ȹ�70Ӳ�;0�e��\�B�����x���1�%;���܁�4Ԥn�����^��n���6z�<��w�R%K���/�ֵ��*l��Gr>9��I8I�19yXSKK�q�`���/�q�ǝg���v��+ny̼ś�P%=����3 *��TV��������}zWa����6�:����9r�v��u9�o ��V(���ے��쒯wsE�U�������� 3{��N.���zi��;��/m�r>����-�9цԢ-O��&�W�c�^���7q1�>�(���^��!�g)~~�<�j�����YEXp��o�>�un�����&��H"'2�GJ*����c�o}�+`f7)���E��ξ��WV��/��� 
�5~S�o��|݃�c�MRڬNc���e�r�/��*��ψ���������mA�)n��p�]+�
_�=��E���k�jh�l��nO��(tW��9cnh8{L�0�:�C
o��Q��:2`�W�d�^ݓ��8Y�ᮞ�e`�%�mv�{�U>�)6��gΜ���e}8nk-r�{9;e�in�րɓ���>$o�s��^��d	pL�j!|@FI_�E���$eF� ~K�,%��B"K������aԂ_���c@���xHa<V�4c����� �+}{��������[�`uE[N�3�8M�"�=5�6o��*���o��7!J.����4>�w8������Sss��m�u]�H��qf��N[v��&�^ۢw�t%@&>9�y6뜥�����O��6���v#^I����T��#k��h;m�-�e��N���!���y���wㄶU�&" �#���̈�P��&~��q w�K-❿d8�\��n����0n����\�ᜨ���\���p-,�VN����S[�<���~��_pv�+�4��e���:�r��F�x��o��m.�m�I���k�y-xQ!�l�w����*g��f�0����-�CG�2?�-�������6��h!�:��| ���wB�y�c�.G�ݿ�P����e��{�ȟ���x.�C��ۻ�Ŏ��GI}��(����9&|��ѱ�)Į�u��m���t~׭�.O�څ������h�Tn�󔁯�F�j�5-v�Bil�����E�'o��4��%��cJk�*�=�@ݱ�Q���5�b�fz�͑��׾xj��0�R��F����r�[���]��p�oӑ����՚����xt۱���V��P<j�
�eJ�Ѿ�Щ����w@���,Yq�T�T؋s )-=qU"����>������:�rY�Ŗ��
�tQiZ���#�c���I x0%$�@ ���Q��^�rx/����Jn�X�Ѱ6��{�Ě�� ��ν�lI�'5�ڠ�*m��*-;�ǵ��������BD'C>��xx���:��Q���-�5���
��ߌVw�Uh;
�����P7u "���t��Z| 5���T��r��1U#c+����]��ŀ�֙�����Q��G��%}�ݏ\��T܎ak��J�������o��m�.�Z���&A7	�-k�&����1lB:.�pP�Օ������^�cgO������i�Rٵ4��e[�q��o�8�$�̾��2����co���.4��JwP�&��}wٻ��n�C�?�H|/WqD���f�'F넉'^��K��ߚ�@�(�r3џ���+9�M����q�«煋��;�����.?m��'\F߿b7}"R��6�E׀��C^��<�eq4ovxv��iH����C��PM��@��x���yzB������*�ae��VóR����®u�xi����.��ͪ�+��~�tQV���Q���zF>��9�y��ύ+6�}���!I�Z*��=Z���S\Io��Ž�֥���Z��ŗǜ�xH(�,h��Z,�6���L�d�=��TU����e�w���=��	G%%J����2��Z����@=999�*6��Y<c�>�'��n��j�Y��?.0�c��j�3�bl3��R���e��r�S��5I4ѓO}��M��et1e�
��ȕI�4�Ȝ���:9��$w&b.�,PQ���'������Rx|��#�� �[�G��E��!8 ��w�<Q�&&&���_N�=z��q�ؕa�݂w�ф3�# <��������y�>diĻ�^��kIl*�j�I�(��ڼy�3.'�^5�?k0�ie��pI*����p��q#�%��<
�B޽����qE�y�+��p��7W�&��[�>`˟�K�tM]��W��uX���CW��N˔�#є�C��o·��>���ͯ��|E�B�sx�/(6y_Zw� �w���Ʊ	o ��J����@T_W��#�~���\q���j��=M��?�)	v��"�b��&V�z@׹�-�@���N��hlR�ք���>�gZ�C����X�D�&�uVT(��9ο�Da��j����*�rO������h3��6��;s����w�8w�Ū̡ՠ���#��W7�5�D�"�U�����Es����X/����L�lC����6��?����Z��h�"����cI��E�"%�PS!����JYCҐ"I��LL�d�(f&�I�L��������=����5���6��s�����{��֥����=�H}�
��X�9/H�c�Ќ���X�
���:yg2����TeM2 ����]���S���T�,Ղ�]��M\�6���Me���X��s>�N�Y48�������W`i6���*b�>�g�$�իW�4L��8jXέ:�1R3J��"���CL�ID���[�z�a[�x�V�x@y��j8�t75��٬Ȱ_�N����G��1s���lmuuC�@ \�uZ~��HAS�r�q�i_i�K�/��8v��W'�GG�LI{:6{�ѵX����~6r�J���̞G�,�S�Ģ�	M���H<<h�*/'��]��������s�<<�=�Ōv��ݮ��^��v=�嫹ZBJve�if9t�C�T���.���t�����ڇ���]sc�:=2������ʿ�f剗����)K�Or-Mj�䂞xL��oow��.�<��J����eVcB��T��*=�hB���C�V�����=�CM�fSD�_NJ��n�j�op�Ӣa��Q�"�m@C��/�v�J�_� d� UO4i�85�5>V�A� �g�m����䖼wwŬ�䅺7�kF��5*���9@�]ųK�8���r��!W׫�bb3�ݗ��Uߨ���`!FJ��X����=r��$�U��1NU��ï׬9-�@?������a����I��ɟ@@��Iu �O�J �F�~b)����{fk�^��"����� ;+qڊAoUӛ�&B�g��+ct*�q�w[n���.𥛫�&x�< ^9��9̢���]������t�l���n}�8�h��s��CiՈV��%a͈�/[e/���9��tL��K/��P�ʢ򀠅�f�m�m
�H�p����[C$��}�:s��KVf����Mh&��c\������:z�hS�
��	n4���_�v�ӻ	��~44׊���j�=��V�z�J1�
��� iD��4�,�V��V�z�<v�)�K7�����F�*��7���c�-���M
Ǔ����(K�mxj��Gu�3� �f)^�e}���F�^�]2��Ke�g���B��Dk�Cmګ��#��Q'�=s��i�Y�h��w>b$9J�#�.,���8�Ǒf��B̊0�"�1+]ă��4BU6�t\���b7l���a��|;�Z��:Ds�zM?"i����#�m�Lz�y���}k�+�E��
r(`S������#�-��ہ��q�2f̵bBІ)� �̸LG��GFP~�=?�pu��j����a� ��W�;�!���z�	ү&���{������C�QR=�]�X���^���5� 2M|-Q���e�TGS)�Vg��Aظ~��}Ĉ+������-�c���˙t�f�,kL��ʵ̱�6y��?Bbv����GY߾�j����nZ�f@��}=��Ͻ	�zFb�ɢ�x\�������~l�g�~�������6!o��	����;��`f2���6�^����mR�#��Z|N��Ɇ����O�V���ܞu�F4���#_��G���D�B�q؟�ɛ.��7X7\��DOx��G޹_J��>̻�"b�R���\D?�M�4���9�?���^��RY:7�S/T���Ѣ�K!����)�+��H���߯v��B�
�Ŝ��)[P=Aдx擘�j�����[Ue������<f�g]��W�tH�%f�o�}iՍ&�|{�;��Kx��%��Ӕ2>�ۂ�����ĂD<OJek}
��1g�*^u��U;D$& N9>
5sƿa��$4��f=j�7���Z��ƹ��&�v#���j,"�G��̆����4�q���\���y��N��ӯ��X���ǋ�Ta���B��'�$[�N)�68xkЯɌ�\�]p�>��P�9��б5��Pd��a���=ڎ�&���"O�u;F��K���a/�9��$���/G/�f�n*)�ŕVˊ}�E��@�L��[��ľ�8�)����)�P��"�*Yqyl$@^��Ԃ�@u)����ɰ]��_4�E5�(~ͫ^@��jKs|V��l��jR�qc�ڟ;���6x4i���K�ىY��:���Q�@�������wr}O*2�Z66���M@������iuS��,h5	�	�w��뱧H�×������ϒ�wI���o�CZ3�K7�3^(Ԫ/���0� e��$��ԾֹXL�o��E�d����א 2�[)=�bq�X�z^IQfX&�uN=�#Z�mob�������C��.��3�c����\~��?rgliү;c iHO�Å���,�	���kϓE�a~@�X5�O�lY�.�(���sq�ۯ��ƿ?A4��t��|�ʑ��ʋ�0֫�7c��Ⲵѻx�滗E:�>�ɷ#aV@=�իF,:*��E%����´b,ŀ��7 �m�R�g�/5ڑ��I��G�[W��+W�L������Q �}�U���$B{2ᕇ�������x�=.��_�B�`�fu�h������%O8\ߗr[��{Ys����R����h�-z��E��[#�m
����5�`�(5i��vx|��0� ��X��g�o�G(��8��^�v i���;/�Ib|=�.��_׹0���q�w7JQ�q2���op>�S	#~RZ�%���\!��̳��|ݕ��!�c�G5�?@�e�:�W<�ϲ:Ӵ��p�U�O���e3o1r�T-�x�1�e��X}�T��ٙ�K�D��+h���̒HלK:��GT��߻��Ϙk���@gh��gdSm�U�B���a�!����ҢZ�[����:=�:�(I	�Vב�~���^��P���H"|����N�H�g��J��e���r�v�?5&���[-c��3O�_.G�?[��T�;nU��_6�pę�ݚ>�Xo�ܻ�CY��1ڤ��G���!=���́�Aʪ���Bm��;�����&/;�n��W0/p���&q�(Ȑptf��;�Ȝ176m�7���5c �Z��i�˖��YEfW��=_��y�Vm�S1���JvCz�Q�Rй��@`I�dP�)/K��rhiSss"l_%[�߇��6!�D��rx_%��J23�v��٢�Ǯ Byj�7��C�����ۀ!:r�ht+��r���2rx�=*�&7���*����bV�+?�(zdO ���jJ�#-%9�������b�)t�Q=F���uy<���C��#�Jgq��!�� �h��+�Z[��ȉ�-���8N�[u#u��A��N`�d���߽�!��g���muJ8�z�pְ�iKXl��y,��[�7�k��x"�����C�1��x���Uӑ� ��́��'�C�AT�\/�����b��-�YR��\�vlх ��#�IU:>����k ��9<��ʡ�3ԦY����^��a�Z���%��e������`���ʯBy�%S@h�d�b�G����	�iZ� aS{-�r"�-^���K��0Z�q��6!�h���7�ᗗ{5ěoT����Gd�_�����f��G��#��w�XI�!kW.A,���~��b���y�V��Y����w�a�g��v�;#�&4�e'p��]@/�.��	8a�;.�M�<K����(`K#I���I�1!ku�H@���߭���Kû�}�.�m\v<i��َb���SH��H�!�`��!ݥ[$)�k;8��ꃭ�r<.���E�NȉqYmN�+�x!">�U�j+.�}7����b}5����y�����l���ϡ_�ɏ�B�鎯VS@��tw㯥�z���TR��Aj���vh����Pql�t��B��ҹ�&H((��R�W2�R����98�owE��w�dԵ�@���h�b��E����ں���Z �����N�����W��Ș����L�BF"A�0j�v~2R֯�;������+�c�����|& ��CķY*���f_���/G�Q��J��1oJ�$P����ש����)b��� �z2u�~t׭�rk����U���_)V`:�#���%�(#5���'Hպ^g�?�y�v�R���o_8��b��3{ϼ�'�տ�'�L(���#[<�i�G�(\Ucj�J��Z�;���՜�v[�jƫ�?z���[R-X̀���l�)y�tV�j��,��
�Y��Ԫ��N1V>��9\�6@�����Z�
�;HF7�5T�q^���6^�ϙ�遂֟Z7���-�Q&J�+����K�w���8�X��}�T�?���tw���OĔ�����ϔ��*�./��T�v�t��z�tl��n���;Cb�]��[}YR\wC��*V���1ƯJ���r+mΰ6��n�������h$�z*YՄ���ܩڵORX.�'�V�?5l�
~aƫ�.����k)�L�˻���F	1k��=ǌ�i���SQHd��T��Ș��e_o&v����ŝ�M�N�-V*�[�=t��]�w�ZL�i��$�U��D��؉���S6�
��ߍ��+v������vK��i�VP4� �q��7u3�ƻ��l�����䞬�B�bp�k�˓�����K.<񖖒]-(]�U_��TavD}��|����aj��~�Ѻ�	�?�����N%�n�N̺x��>iw8��{���F�9�p�c�22V���t�'�'��H�����Y.�ŋj���v����{?��	�7������$E�S�-��嶺^�M�M�
"�#��i֣�]��Q\���B*����u�ۥ��U���Ք>�(��!�T���WR�z�a:��B
�
w�u1w���`�	�t�	��(�"E�&���m&���;�#Υ$1���L,��*&F����ݼ�rs=˺�!�����y2�-�-0�mw�?����uA��<�?�4���]pz��I��y'�1~���y�s����ս�a�%{=1t�Bb!8Y��#�n��
h�g��GO,_d��y�+;)�X��6\�����O+�8� ������%��>���*�,��J�e��g�Nt\U����V+��r8�qx~���߶g��,��b��{t�W�NɄ =,3�~��[+�Z�j�)&�9�2G ��ˬKA�����	={%�]G�?,�rM���7�P*��^���?u{��형q��T���s�ݾ�
��Q&�;|���A�̨p0�f�0�mB����x7<6�� R���(�3D�~�����B�ѣV��j�~8�����B��,�Y��b���x/�w6������i ��KM#��бF��L/S\u��W�s�*B@U�����r�i��`	%�& IK��2vY5������չ �/*%F���`����̜u���	
.�r�R���hK���+T(:� �S�����||+���NLU�9F+d
1���.�W�%߮��������%�!t���fAS-�q�|������J&-�N;�m)~[,�o�^��5{��pjD:�р�>]��~��3�����¶<y���H���J�\>)�(��r��OT�v�a��L-�jOv���'��3��ź{�'�wDsk ����k����u�K�3�l�y����V,���J�d���Ƶ��W7Z�`�5�������0-8�M��܆�S��>3$�v+�W���$��O�3\�t��������[����~
ǻ��W���y�[�k�b�oɾ�d��nh�;٫ =Q�u"сou��+�t��f��J���P ��.8k���nu������^A�8>X�z�ńr�����h���_�{_̼�cb>!~]�oG4-��%�'Dq��1P� �5#�Jh5�!�9���==lAȔ�i��� �z[�,��Ru��_�ɻ�p�3�c��f�\O]!,o�e_,H�8HC��}=�eI���0��|�Nu�1T)���ӭm��IQ��۽d_��h
ba8�a�D��dlh�� ���R$;��5�d�e�:h�Z?�-�˼�0�a����9m$�w�c���k���+��̓hM���?�D&ֽ�M{{��}�u��c���['jÖ1��?�������
�Q�{�����6,�&|{���3Ͻ���:Tҩ��Ru)�}�����i�R�L��<Sr?{*�35�'~o��g��p6<�����& ֛�JN@�)�_�t�Y?��>��9B	i�#4��~�j@L���R�g°q�N���e��,$hfv�`k�POЗ+|�>z�:�X�b�jg���(�f�8+q�����f�Ǵt��4�)��Lc�9�i�ًS�zN�Zr2w���|���v�����r��[ ��o�R�v[џq��ϊ>��R\Vq�נ��Ƀ�yv�,���$@�AP���������:�_+<�S�^oŋ�m�}R���7g$%��"u��7?uV���s�B�^7�`M0�]��B��I�{�A�k����?^�[�`�B)��^.�=g��x�?��"`���n鬼0�p�ú�*Z;�B���%8[`12��T?*�fǷu�l@�3v��5��6-���A��(�'�bJoV�b�ё f��;����T��a)[JW� ���ȳ�+3�
�BUW'���.��vo���\,@㽉�&۳r���ߞ.�����ޏ�������}�����Ѽ)���<N�I�R�a����ODb�Qx۩��e��b���%�nbCNu+������=8;,��s�T��3�M쮆�fc�7�()Q�������&�LdT�v@��6�WN�/gT@O �F��*�L'ԉ{���M��]�ő�{�Q�'��D��9v�K?��J*�_�d�B�s)��L����X|�N]j��\�c�P�/���ć$?�~��$A4�Dw�ϯ;��� �J���;^u�Eפ���5�X�;�	M��`l�*$PW�ށ�)r���ѣ�٬���
V�@ >D�J,<�	�:*���@6��f��o�Y�fo���,W6��Y��i�z2��z�q����3����E�">��<�03�ڦ�HmhQwE�;�>*t)�w:WD��:�ǧ��g��?�y�y��~���� 6.�����~�Tk��(J�*���ʧZ�Z6S%M���eB*	�Tq[�?ҁ���r��Xቬ��-7�d"&�qo"���=���**�O��su��ź}�z�B�����cCo�����Q��9#��������:��M|<=e�R�t%&ȇ[����W������K}W#�J( ���;�O�?�!��ղ���1@3goS�6�e��;kW�} �I��ZЩ8�?� ��V}�|�R?�(U�I�+�t�:'a�AiV�^i�ڏ�PIg�cjn-��/VWڥK�ﬥ��o&6����$���t�<e~�^a
��ct0���k�h#P'�%��|�h����GN������_,2�{��
eK�
��$_�n_l�{�f�ы��+��t�cg�m��s�%{��"�1���=�~+o7�s��G �!�D�g,]�{X������6k����O12�Զ~���ș}~; �ӄ�������� ��t�?h���� �Ж~9oxf��Y��?�f߃�w���s��_"��FJ(F~�Α=w}`ک6��P���©�����a �#{:�?t�D|�r��q}�s ���:�����y�B"���.x��zdb�$`� �B�*]�mj~�����ν��Łe�{�kQ�]L�����z����CtP(��Qh��;#!o�������ڝ~w��������h�lP��]��/3L�� ��ܧ��ԹS�]Z|.E�6��a~�e�����]�ɋ䲣�B?]���8�+vbJ�Gݿ?	�� ���,$	9vK��6N����b���������]5��^M����
�����@����ҝ5H`q5#�^eXؾ	���Ӥ�Ö&e�un�����j��4���),u=W�.x��o��{�k0h�(�� mH!1�֕��Y�J̐�Ke�j�|0o���B�
<��e�'�e+v#�&�H�E1�Hd�Lt{����b�vHe�q����N�j��wR���k�LXMB�h'��N13���?��=M�V� �v��0���z^�
��%�ˡ�h_tힸ�Y%˟��Ɏ:��1�A��!P:R������8�C�M3v��y6�駚��8��n�!�U���Hc�ͥ��Z��À�C
�?��w�Ub�z���#O����G�٫��{���i-E�]�K�`NO�} ��T�����=�~��q���e|y
�%����z"ӟ�!#wBO}��-�ȤIcJ��!���S ���b5r��ߍ��Hg��\�x���!=\��4#z�5��b%';�'Ǵ���:���#@�9{ŻC�q�p��lzk���d�����Ǎ���P�ݧʾ:�܋C{.!Ĩ�g��/���8�|nS��u�*� е�;2��X�+���	g>u��49Y�*ž ?l5��e.>��t�3H�쫅�_����m��E���M�S�7{asQ��&ߍ�{͛���.+y
墸���׻��)����=V@�kӉ���ׇ� �}�� f'�7�ҵ?:|G�4��U��?���\A�)�����;����u�.��V�{}DFZ;�*ҋ����w{Y�P#���>���9��5�%�;�(ܷؐ��A����cQ�t�M�?ia� ��Kf��ݰg�ٹ}���S��-p��)��t�������ϳ��X��;���k�E~Ї�1�'�N�e��J�?����v�y�}��Ld>�����h�V뉺��pq����|i�Ap�f����Ɋ[�������jL@�vx�6�t0��m<���yi�־H�Q���7�($�Q����NqT"�l��HW���� ��3������|��ļ��B�2��R������_�X�����y���(�j`Oɼu�D�6ᧁU�����פ"�� L��X�B}�R�x՟ZD�nF�Υ���y�i?~1�Ke�n�� IR�]�&5����7`Ϗ��2�����^�^��X]��>���gR�@��.���:��J�� 8=-GVE�^n�L�']��4��T'|
�?����*�	pf��ҧ��~��(�ݏ3����+��=��gjbsL�o���ǔH���Tzu�V9��XIL��a��*|��D��[�9��m�_<N�cyk"����.�3���zw�d�7�d��s#�Z�J��i�`E8H,a�c�*|���h����?5>��-���@l��yp����f�~���d�vM�F��P���xK��luM�{9yyViii�����3�&��չ���Dl����ڹ&|��=cI/����j�
��'|~O�gn��6��,�Wa=�֢P���㕋Y8�H���}����fJ���b�m�?�Q�Ҙ�����?s�u�?���Q�¡P��[�8����`�I��nI�������֔ %Z��T����������t���ks���<��lh���ˋ��.�8B���z��Ƙ��w�����V'����F�]��(��1%�̺��S����,�o���������7yҼW0[|_�������G)�,7_j~���N�)��&<"b����ŭ����)$��#b�Eі����o�pО�7o
�h�!|�*#ث{�^��xXg6*@�_	�_,�2��p>
�j��҇r����hK��#�󌠬��R$���
���dJ�&~�5�~\�6pB�xu�')�os�@���Q�3f��a4k=k��g��}��=�5k�a�Lr^�<�G5`Ệ�_�8'�lW.�&�+LYP#(//���NrPbX��L���\��v#XL�1��CU�t���2�$:>����u��so��0�#:J+�Z�)���f�v�	�U�Q(���f��پi�Ol-����:����.���~����n����=���4Ow^C�����8P]�a��^��[^��6�ΘzW^�յ4e>+{�釄ͦ08ǒ���&�Q�F �p�H-9�UWg�f7؍�纠��6���)��lzb��+�"C�-�Ո�CO��.#�zH����y�����$HS��982C��TE�z~��$�%�C�e�Cʢ7��ق�?��tDy��>j� �l�j龢^,G��{tx�o�{m�s�()KvVz�	|n�#�@><N
j���V�c�׼�<=N�er|}}����l��R��7G�g߿��{�=���������B]��>ޛRZn�ꄽ����ɦfA�vN�(��/��1�ii�y��yBI~Sv�˔��Y#v��fk�xi�rqmq�u�9/�#?���Kv�f�|��3)oҋYG��i�<�����oF�����٩�P^N�Uϭ�w��ę���졔n)�3��J��q�$ڍ�[ݛb>U`1���C�T!p,2X8nC�S@UG�:���d�n�����_C�6zN�[5�)�S�-]���#�L�`R���x���~$�������M��%og�6�ۍ#�r�R�?fpXuuu��hqU�l?�7�����,��5��7<�w�c�kf���Q���<�Ѽ��_�M���0d�/Pg]S_��H!��&���#ؽ���>xLfx��X�U'�zW3E�O�}�����Rm��
߁u?��������]�a�GD`��\w�&o�&W�&��o���p&X���#�!E�~uڶ7�롼���>)K������"y��G���*.l'}mB���������a%������87S�;��F��Gy*)���0)����9��7d�rI(FY�DP��3v6}����!��\�?���L/Yo�M\�
��p��O�
�N=6}�^z4�KKy���\��Ƒst&F�V]�;""����TL�����%a%)�¥[kki	�{�aq��8	�=�,���H9�߽��� �u٠�*{Jo)°! �]{���#@�v����	<�@�s�*(�od�CtA�\?���������Fy��sUՑ����@�ViIpvn��lGR��&2�� d��	AgB*JTN�i�S2<<�ǔ��KQa`��J�J�PD�A��%�m�/jiIx��-�ۼ}�G!]^NΈ¦{� ��^N��D�a��<n^|d���RW#�&]W@Mz�����w����F���vy�y�=��2��Mʏ�<�qk����\B�D��-_+�9D����DAsCV������UC�To�eX��R	��y70���Vu!��g�����۫ et1�����Á���@$�37���6�O�Shy
:��
�N|��W�vCV-D���R��t��vf&ZF�XIiV�������:?�$,�����dO>s�^�ܼK��G="<�c<�Qذ�������W��|-�vv�$�׉��Y�2���X�i��	!����{�m�kx����@zq<ye��)�b��(wg�O�&W�Z����>nv��#~7~b�ؒ�^F����;�{��0Û}���݃���~�^^^^`v:�C�p��<R�������E0Uy�jj�1�zd�Ei�Ztϙ��c${qZ#Ō\p�kz�����Ҝ�}b1����Bʵ��2�)��3�3*�E����������1��vY�2T ��M[d�^��~�����6)P4g$|?�^M����6��X�}�䱨4A`Is��\I��ϲt�4pU��5
<����1@�J\��8�⋄۲Έs�ۍ��N`!W��I+����t�#N�T�$�]Ҷ����=*����1��J[M�E�D� k����ҫ=���E����� ҁ������O��5T��
������MAx�H�s@_���͛�
��ԗyIs9�������m�s�k7��ͬ��r��J�9f91�Y%i)sH��	�[C]�L��� m���[�jy�#YF�|"=�W0X�u���z}��}mч�OY��I2�\�����"�Ifp��P�͎��������0)i%��eA�ǡ|=��Ip*����4��?��p��{oZ�q]��x3vX�סFΩ�SRƟK
^T�x���Р��R�Ē�>Է�o�aI�t��&7yIw���'o:h�B�W������������j�\�۔V-�rwp��o/�&�i�5�JAeef�k*Q?����iao�9�d��W�&�d�����m��d�&��2J�����۷�պJ����V�H��������� �x46�[%n�L��RU����\��a����L�� �PFr6����wUP����ѹ�����?:w
,�*���߷~	��KG_�]�'.2g׋��-%���,`��03��逄uqQbi�3Z5_4��G��y�
��g2�d����#�ы�Ǻ�=����!,9� hj����0�:,�=��f��2@���8k�s<�ܮ�0ނ�rkk���Ѣ��c[�P~����G{y��_.�N��������$��v,LV+�����FQ`��q�";���(�!.���;�|�C�lemK=��;;���d��<�]�2>�����_YXX�e�x���h_ld�[��������K�f@I
yI/
�5\�O P;w! �e�Ka�cxj����i���lҬ�p���0�p8\���Z��=��.�eغ&�o�>1 ,<<�+�Zҕ���1�ض���%s�����P9DpM�E�&u�3����PC!r���%/Ǿ�6`��8f¿�ͦ �+@�H�� ii�eO��v�I���ب6�{�s> �I�����Z�y�Hr���jcAɅ��2&Zu;xT�Oj��A���^5>g����`R�ֹGK�uu�@����F��s`C^� �%�VU{���򤏥����MnI?=�<'V���6�3���Gq�RfQ��U��Ǜ�W0�H��顰�0`��Qc�w�Vb���u�[t1���ȶ{3δ��J~�=���t�)
�jqZ�8*.���r?�-��F^^�Ƅ�GL��D�XS�#�>c�x���NN����Q�^�U�[�����3��h�g/�g��c��"��~䦽2�t�&���"@s�Fq?��L�Bs�.�)�ޯ�W@K/R�����P�(��a�\&3&�B��x�BN�O!3�S��$��$g�g��/Nkik���Z:�bL��g%��Z�﯊l��h�XF��R��f��w`�ųYLI���|㛪3�փ�Kva���R�)|MSKn��w�,Y3����c��Մ<�EXY��K�-<��ħi)��@,��Ot���r1�71eп""XN&�y����o:t0	����z��:��t ��ny9��6����?��]A�aSy=�؋W��2�>�垀Z�NMV�[U���LP�!�miqGg��Հl;Z ?�֮.--��b+++s���;o^!��P��1�
r��~v@Jgz��H��8���a������|<E�O�v���k����*���8썰���;)����/����UU	��Z�����r�3�$������-��d�k��J��G�$a�G���*u��/݁Tx�,~G�S���/ڦ�n��җ���O:]��c��(��,��>�奼�y�ɾ���*h �$�Y�e7I@�u��j#9:-BBB>���,�:"-J�
���e��is�Z�O���]�^[6�rsA��\��&�_�'�,��s���O���ԥ7
�><�M�c ��|2@��A��VP?��|�55�@ q<P���q��2��'#9���B;
(sW��I��P���t@h����s%����aP��2OvxPc�vmwװ[C*�I>�/;!�?�;���Y-��xx6qEaS$����54XQ<�,)@�feyk^�AT54$��=(:�K�+ �$#k�Ϋ��mdl�������i�" �j�4��������/�s�ߐ;�V��N��5O� ϯ00�����y�`Ag��0.߽��܃� /�i���77��l�~Ɋ�����~.�-����@�p�����3�����! �T}�f��~��^��]�!l.C����,�wK�Q�������!�lf���W~<Y��d@0�u��@�U�p��=<3�6 ?Z��.K� \�?7���g���)�����|?T�W�y,t{�$mi~#rUvF\˷���#�=��(#C���3���D��QYH�I?`S���P��誙M�,H%phf�ثcD?jR{Y�����6@�ϴ[�F�m7������G�o j��*0R�SSr�BM����Gt���~~4�>N�GIH�%^�0���m@$�� J�P!	�rKKB^�f }222�����ʥi��`F�)~߀et��} �=f���lj�Xw��C)��ko:��*����tM+�{�z��	����{U�;~�0�:ϓ&hhX�|sG��[��]j��&#L��q2%��f~?v��n�^nW��k�6�2��Ky�f��}b�~���3����5Y9#fzw�5@s����g�}!�y[��C>��в=fi�jj*
��ǿe��|��彿G3��(�&ć�*�.�E� ���o��k���G�>������S)��`+%�J����8��F#:��f�Kyϖ�4ϖƱyv�@t�&��������:4�ݶ,c������V��d�8�7�I�PZ���n?H�Ibxg�`��<罓���f��k�[6Af��f�a>H�����7��B>�{*w����Y*sC��dH����J�qSj@�qk��gE;=�1�,�ТV�($�¶K��Lxi>)Jc¤���w)�;�S�0!�֚���oY��}?��V��=�݋<(�`��+U��A6
�MG�ab�U���4����xJ5�d��4��3W��~����E����N��X��������\Z��
Cɝ;?l��>��^w J�,���:��孕y:���aBO�l� h�4d1��G���Pϭ4����tj^�+�W�Ɲ��,8.(���#����ʢ,�'�r���n/O�h�4��Ǻ���F!1�b�ė�g�_.�BD���?�	@JG��}3�#67��3���C�uo LhqPV�BNN�����hi�����H��
����*����kg�Q����6�֛���Yr��(�钣>,?�:!50�ڐ�4�1�ES���<ξs���{�VvSÖ=dp(�:�:������ӝ�8ˬ�!})ː�7��h��ԫSԓGr���c�-�I�����o�~Zҧ��֫��@=���C�X��fxh��<N���  ��#[xm� IGԒ�(3/b�� q���5���Jh�|���2d ��f�(�}���S��'Y��Ӌe��}��=As��w���Xw
#��/�Qcccp(�� P _6{D%�Q��Yba�&���X�O�3H������{��H��7J�Ez�
S�vC�r�5�ح�{P(,h1A��G�d���ϡ���	�؊��N5�ޣb*�\
��D����X�NW�oӈS��)OdT(�|ρe�ّϦ�غp�v���e@>Y���� *�fˀ%>`Q��#B�G���03-,,�?ⷧ��]$�6gط��ny���l�Ps)�S��E�8��Qm�@�E�>��oM
=f�d.�������3aXG�	�֮}
࿹��͢��G&ES�����ɓ���mX�!�ʉҰբrgM*0��Q��8!{ďf	����o�	h˰X���M�+��{�K�U����E~�F&�v,H�m�����e7o:��=��z���8�{0"�%�r>Mc�X�9�Z���:AKS���<9���YC�)K��۷�\��<�?�HE/t��M�t6�rU�^/9E���铿��J�E��b���> ��,kk�e�2K����q�.b2c�
���ҏ(	�x�Y����xY��|���:���t�
O��� $� ڙ��?<H��{�A���+�ol|�#l,K��q��(�M55�!��X��+�g��Dg&��|�����tz����~�;b"I��7o�s�������I��#�֌:�
H>Es�>��i�) �ȴ!�u9_J&[�S� ja�p���NlqB�jVנ2[�D90��b�F�e����n��yf��y�_q @5yʰ���\�G��Vn���ex��y�IZZZE��:��̯�����3�Zɴ�8�Eշ�|�W��$ ��yl�D���� 7{&�X��J���/�}��Ԭ�w�y�|�g��G_{oe{�;���b��g	#�:F��+�Y:��h�	�P3�Uw����H�I�Ll�$g'�NU�z=�4Ap�$�pxbȨ�J��V����ɓG�(�!��{>�Ds�!���YiG�a����o� �{ࢬs�Ds%',�n���W[D���)�(�_a��t��9|ԅ�f��{�E�$E.�<e����5'�g�f�O܊ᭋMs�=�Q&s��ƽ��)���u'C������7�)�?r���C.�Գ�b�gͯ���xg�؛��I���W�8��kW�y��ޚgsm��c+�K�]����ߺ�k�_����3�fF������Z���M�"�����j��>M1���n7�L/�^��5!4��	UZ�1R�_g��eETN����?�ҾM���|^˖���ՆU�z��Q�Y��U�*�]KS��b�ɫk�-��eP̂���y{n#Y�q̈́un�=���̯�v�����`�e�0�`�V଩}�ڶ2m��wʤ�k{�r�p�[\��s��N��S��-H�*Ƞ�5Ӌ%���׳>b�L} D�F�E�!N���38��?Z}���e�8?��~r�gfDs�Ϟ���Q�δك�K����K2��&ά��k;|U1K�����V�G��#�+����p��'o�ǂ��Ӻe$�G����n����xOB��X�
m����mB�c==�\gn=���?,��5��8~�u�1&�����$��$��#��6�u�6JL�^T�cg=q=k߲�$�V��KH���>�����Qٳ��r$�<����vq�����*iA�q�V��m��{,����l[d,��Z�q�h���na�#@�#޲_��Fs��O�Z�����<3%[�����2u͏2���w����6&�~��8e¯�0��~�z)�D���oM,Moi��M[]���W[�6|T{�̋vXs�m-������;�֛�����-Z׬BW�]z\|��2-1�=-��~?�,|d��E�݊���5�iS�`�e�exU ��~v�����xO|x���F���F�ZQ�l�7ُ���L��\3���Gs��Pٳ�Nt�;lP���6�
!�kx/����e���aC���G�e��~C��5%Y�O9�W5�"����Ƒ��ä��n�r�n��cͼD�x�qrw��y�F��[qqqzL6�0���l��+X���j�G1�Z�M�	��yX�����l�ph5Y�� �%D�P+!�Z+���5��@�b[Sa{^C����:��=�û��m�H�</��yգ�h�P'%+��i��G���-oUe�T����?���E[���V �+b=�%�`5}᦭ ��V���V���]J!�3���U�����(�4o��eJj�k�~CCHƷNfYD姢� ���C�)�3���;h���!Є��)��|?���Q�f�d[ۜ
w�XaV�q�zd���.�@��,x��8+�
��E�G|��M�m��1	pC V�*�XO*������5).�G@^!�~47�00�ֻ1��R^���e*���F��i`��g�)��z�D:n�=�d��ràL+�h��e�	��%ߖ�Z���|��vͷ��ֽR����Z�c��C[�hn~��pF��)S�I�u/����!�$E�pQE;0��"R������i�-���)'g�+s�?u(�'F2%.��W��H�5�	C��"N�> u1.�,���pc�Tj$��'���4�ܛ�5�{����:|��e|�����$�N���l��)���
�G<~���3��ɳ/"_�gɔ/H$Wm]ʻ��N0��ch��W`>�I@�VI�s�eU�{c����b�>�O�?���9>�b�T�fH h97G*;�G2QO�z�]nU����$`�{k�T~���	w�*i�&�YvXS.�|��`+�,\jz�'`{��F�?RHgTm
S2$�(U�M��6G4������ !����C�<�A�q��!����k�f��,�E��m�� K ��:pYb_�e@�E���H$Y�ٳ�0ؑJ�5V�0`��8�3j����[A��`��ݰh.X���j9�c�ݤhġ�.�nQ�*�3*V��s�<�:`�����J�۽�H�<$m���.﨡UlJ��,�M��c;�w�aqD��w��?��2�n:å��Wz��/�$5w�|
UUmL�X�y���ȴK��u�8�>l��8j�����D����UAo�zo��{;�bn�sr.�&3s��h�cʃ�h���-vBȉ�%.����>Xt��3Hh�W��h;w�2����57�KKƸ(u���C.�Dp�D������\ ���.�:������mUW��e{W��86�Ͳ�ƣu���Ç\�8pIop�=Մyb�]@�/���a=+���g���c��9�m�:�.f?a%O&~�J�1_�A����0#%�<_Q�TD�`cv�����?�y��~;^~�3� f?{)��=$W/�گy�6��4�D�H��յ)�/��EΟ���P-�>`ViE��?�ѳJlz�E)�����d��5I��Qu%I���Ӄ��y��7D�'2]�����Y��$θ�v�t{5�:5]�q��8A���W7��W?-�:����,7��cr�w�	F8����^`U*v�=���6��&�lN����I�7�~|=�Co��b�=ɢ$���X�Cj�m
b�<p358D*�loq�)�0������{V���Bw����2���Ϸq8��?9p,�U�1W/��^�\W��,����ph�^(�mՇ�B�� �,�������j;d3��3|��`7�- Y
��_ң�nF�"�y6z�o�����\��̞��a�/m����x)�*�lZZ&�1�]/RYc����JM�1�_H *�
�����p�V��!�w[,�$��7�6f���}\�$��nm܏M���� 'Ty�w��z��PRU�c��\�1��_TE�9ݕ�]�*��"t{�wV��I1Ͼ��s��x��!q"ab�l,�����y�y�:�)�MGX �d=���9���GL4Ͷ0Nf�)	� �F��8��\�$D��ǜ��|Sڞ��/BVW��}����К4������1��BA`K�/��.����񉯎�P?���JYv��qY���m�  �.ِc��)&��.�9`�a�w@8�Q �455�l�e�{�8ɛl�G�=�ѷb�c}��UH�C�,/{�����%v�g���	ӵ����Z��R��#�Ϸ�08������$�Ve	�!ч� �V��Z���g{�7���eSkTTT��A�G�0�4���晫�E�^��Kp���1!G�h6
I~��%��h�7ڿ�y-�"�	w��+�"�δS~c�hQ�
�U��N�h�[m~�}�>Y<�T2q]`�5�w��<ߗ�"�
Ɉ�	�	i�K��)2/wQu72r,�u6�ؑ����{?��1�޽�K)��y�o2��'�^��jn|���4H G��w��ق@��=��[Vv`�벇 �?=R|���,�P����2��E������s��P���C��D7�%�v^�1'��	a�$�F��rz]�hŅ@!ۃy��� ����{Ҁ'�`Dyﲝ����e��@~U��Mw�� �P�����j��{a83�|�ѻ�?70�.]�Q���_����'[��V��XZ����[	��t�ӏ�_��ǹ���)�f/c��y~ȅ�D�IG+�E��W�*��(+a�q""R6���\������)'��"��u���� k�����mm�J[�Bk��Vq1E�Xe([V�8^�Be(B���"RK-2#������D�����$����_W������y����8�<�g�Dݬ�p��L$�`Y<i��͹�3�e��ĺ�-uJ���<aV=���0���M��t&��V�c�w����mS�-���k��<�=���^@���WWR��\o�V�ٍr�6�R���ե���\[���6��!m!��ORZ�s4�C�o�o㒙��זe�nx|FBBB�����P�D�Ċ���|e���[F�IS0!Y�����z;r+0g�~=w���q���������P_�����
D0�X�J���ӠJIBJ"3���e#�Jj��Y�N������o���Nq-�QN"���A�?�&,��C�@����v����ɿ���#��M�b�����W�G�Z�����R�-5^�|��gC��:��X�ՙ{	�&�S9�zmɵT�2��p��}��J���:�\}���ŵ�:::�ݲ�տ���,�����8��	c[�>�{E��)�À�M>RC*5Jx�}v'��``��Z�#��j������A}�A�$�S��\4�l0��p�C���64D��fgg���CN���8�訹�[)`Ƥ��GF�\��p���"i4Cہ�؋�g<H���+��S�i �����M� ���d�C�_'B (h +:��hT�.�	8�ch�!��F^2�*LiW�!t�:?������T%�) 3�Q�C�K�B�p�?�b晝PXB�~�l֊��-|���i��03�\�s0�>��X�8����
�un�unc�H�������u���A��������Om6�Ѕُ�����\b!��>d��jF3c����M��=�L���$���"1�$��r��Z(��TN+�L�+�h-GȵO�������.g�8L���4�%��s�廂�k���-�vSB�8�Ȫ̐k���!������@Y��D8�d�r�`�y�������g���� ��%;i��Ƚ[0�J�끈	1�MTO�o(�Y�O��!q4���'8J�5�H%�7��F����)8d�� 2[�´h� T��Ӈݒ���Y`�lha������VF���0�z��t�Z����n4�����{3����K4�U`)�c��Y#�^j���/��}�Ơ��{�w�w,H�F{�,���a���c!���>���Q��GG�������Pi�.�|/&"t���k(����1:��۪�'�_����(��A��\>Og�4�"�8��ԟ7�'z��؂$��\4"R+\�����hT���"�p��|�;�q�G��X���KkGIk���i�$*�	j�n�W�� ��B�
���ә�	U�����W�l<�"�;d�)�a����Γ��m�ܱ�o�W�cAr*j�k����lnn6.�Q�nf�_��r�߿N������:8L^,��»��Hmx�
��>� �-�0>=�\��;���F5~�v[��nml0=%� 3���3��L��j���]m0O��u*r�#�c����i�����k;�q�� �Ǳ��yi��6<������0;Z��*�9���M=y�����e�i���-@l��Z��`�����D��N��_7ʷ��֤͚��tٱ�����J�k?���o4*P�}�'���]"��H���`ۓ)(��*#7����dca��b�"�>в�(7�Z��l4�����gw��>��qq3�I��v&C���0O�N�+����U����k-[�Z�5�rRg�ʣ�%��Nx�ਙ��kc�b��h=,%��69<6��;'>��ȼ���䲀���P;!�(�� ���T�l� AcŵF��77?�ܻ6���dh]����0M`ֆ���F�[�����öN����n?�\�X��c�6? O�ҙz�£�-�4����<�4�־^Z���A��n�1Vޞ�H��{��Զc|[��t�#�1�[}�z,z���	��z���|l��|�֏��wi�n@-L��<i�>1V�Y� [p��*&�Y]�>����"�/�l�r��q�섄�ڱ�m�sC���|p,+L]�W�h�P�k��h��P�C�����y7��~w4�Re}R�O;��4Q.�S�5bO�{0���*߇��k�L��0�n|��T�DSV����3kIz"����]��'����JP�#m֦��#?��>�J�g]8�8��S坤��,;�	�6�MP�ãO��E��� �2tD�~�HBp���j]m-�� 9�r�Z|���o�,�A;���&A�,fvVQ�L��8�g�a�z�t�t~��@;���Tp���Q���+n]!h�%�joEW��v^�k΂�@�;:9���74�2H�f��~��n�Q5��Dm�����|tUpp�� �Y��U��~��zL�c�� [���Z'yFʒB�~�]>hv&~]X�����7�*����}��Bs	�5�eg��Be���پ�V#y���j���ۇ*	�g���c�r�ǽ9�ǔ,vG@ȂA�wQ2�)���\������PϜ�N8s�Y3���0����������BD��j��D~>����3N�R��u����fײX�q�D���[����N?�D^\�=B�D�ƕe���oE�|���]qtZ+�h�րB�����G��v&�1$8l]5wFy�[�����Ed��T�r��u?y�_�>�����^3���l��ܰ.P�	����j�-� )���)�t��ъRP�=[��N6=C6u�`@�a��ċ��{S�r�\w?�E�	A����X�L�d�؊����<��T����&�H��!�*U��b��0z��|�z�~� k��u<�Mg/iޖSa%�-bs�B���Ձ�d2�3Y��S	`����,���F�:)�Τ�Yw�*Z6%�z,�_�"�ePX.X�H:�����p��4��@C����G}䗀q�(I�N6S��RY*<��>�������Z%K��l ��,0�ԯ��+5~(�V9ಕ�þG�ӽ}}��_�Ǔ�P���V�Mqw��Mbz�� �����O�+��u��N�b�2���x��Č�N��:;��Y5˴Q{�͐�D�$�t"~:�yQ�Q�ה۟_��j:Q�o"0���1���q�a111�બ���k���?�WYk����k1"?�(<���RBy�	�6� �r����N�wӎ�_����_����v���~A�3��(�g����=Lب�wb51���8������	x��<GM��?%�Ǌ�e��A%��,]5��7x����gѝ�&�����(�P*����@��=2����s�z���X�__��ŶHC^?����}�Z 0�ߓ�$%�-	̑�j��h o��:mc��=Lu0pj���cs�������y��~hb���?m��$G�^��`��:���T�_
|����ܶN�	R��t�Gle�B�
�QR{{x�p�LGF�B�sk::~�D{(BZ�O��4��zS�����T�\CK;�
sS��;P��-��Ix@B,E�X<����%$�f�񙗝ᔏ�wb�CP_M.R5�M+M�_���L����!�9�ܞ��~��>����\�%���ч1�D��0�$�_�M���l��zb�r@���;��7�=x�ժ�������|,���mPܚv����P��=����ĵD
��=�_α�E}SS�57غ� ��SAr8��P|3�G�b߼���aG$��?��RR��\���:�@�K��|<OC`3�"|��d�������!\���m4Т��t����C(����g`G�U�fR��0?�F�I��ml�B����5M���}�������"�hKe�^��dk�oGw-[8�
�>����ɕ�_���N(�ƻQ�>�Z�@�37,
�9�������?Cs��zEm����k�L<ܬ�n+�ut��5;4�
�4:��
�"�5!Ԃ柕������*����2�J�>��2y�����f�u���P?_ˬ�����vX��Uu�<����D8∐��� /�+�7g*~�����iT����/���)�6�x���իi�q!-�[h`R�]�6����9s��S��zKk�t�J�N����L�����
(�<�Q���/B\��h�_#y�a�����V����e趽{�Z'���&U�0r�Z�?�^�0�;�*��I�J�Ty�������"u�3�JP�<���E�|�Ǳu~K�З��D6%��κ��>���PU1qV����&��2z�y:l-q-������L$׵�Ŀ��ՒhS7�\577�)ײ�'s�0������c��fh�0������Q�W,�@�M��q�ϝ��I/�m� G!|���H,4��D���$����QPo��4:wD��������y��	��$�Q���X]��H�4��/����3�a5���!�OR��2�Yo���iႈ��*�r��p�`w�m�+n��������7?�cD�:��~�G��o�A�}~T
^C8��w1F�=-!j���7l
�K���V��H��G�C*�:��W�/B9��J�}�Y��-2RWv�R�
�żj��|��%@���N��~��	�C��7�7����7�bWd�O���i������U����"�7��=�W�~?E
��{�02��Yak�/{���<K�У��A��5w���P��qd�[�+ݑֆD�,"�9�,��N1���Ԥ@��1�zĶ ���.��Erq}k'?�x�8�_��d�{�M��m�C���o KN�W���կ�|�i&;��u��)�2I_�	��;2���J4�!�/�Pƫ�����hȳ�q����e���A#�:�xT��p����d���y��@�W(�*�"�/k����h�>��?Dʨ��bJ�T*�0R�y�c�K��E,�J�p7�l��6/�*�-��C}u�U>��N�W��Zg$��rB��)����)}&�{��Q'�ޖd���H���tt������|J'�����^il��}�Fjם�����J�0�U�־�=��Z�Y]M�m@�9�dbu�u�9xZ]U�A�)�A���!?�/�{�[*G^���J�Kk�l�)�	����\�9ad����%���̖_9�KdC��&&\�{?��Z�_O�0ݜ��8��Q�6���ֿ.g��m�UY�zaJ�'��
�V���̬�0,K�����E��-��K;�m���1[%ȅەv��O��!�H(�ђ(��o�b��BY1�r�Z�]m��մ��_p�X�[C�2S�{�Z�s�C�R����Dn~,�8,u���?�:�4�	��b�2j5��|��:�mu�"/������隣8?B���h�����BvE��x"gl�{<��/��Xݝ�+���������E�B`�Gd��սW4��H�_�^�$�Drww'��ǵ��y�
!���
�9u�Si�N�>�͌��%T�`۲�R��k�����|��#o+�(T1w������y�L;-8k��𺃶~���Ed�p��ѽQ�=7���L����Sc���	���~&':�q%��]�w��g��e�Q������0䵛U�W �T����a�K�h���`qY�I�=Uџ�o�<
-"�yf�ͮ�B����B+
�<�{#u�uA��F�a:.)����D^�[�B(�mV��|~D{4uMO�%�g�ǭT��T����\zyo��N�ߪ������!�x=�B���-��0���'�ۦ�5���'JVM���`�p�v_�Hl����hhh0�%���m t�(n!�XE�Y�^�zKQ�M���S�._�~�,z�AdT���&1�az~d��ߝV^���������X�@C;�7��\,�����3<Q��Oi�ܶ> �;�.x��a�~9ڄD?��z>�U{�t��in���ߦ7�����V��f�.�8�yv�Y&�dQT{Z����C�Z]�8q-��X!7�E�!�
�4��N�5�����D���5Jb��\i��'6zN�K�6�;5=��\�޼l]�����޾x�,wT>/�ez3s�as���ZZz�����Sn����\��c5���r���0�Z�*�NT�h*.T*��Hԃ��w��[�e��Z�%Q��hB��ʠ���������-(^Ն/��Rs���~�D���-��a�&�~8�*��[��#Ճ���ric��k��3������ @�B�̺:�2�H6Y�`(���T3$Y���'����/��*�hn7}o0���_T���چ1�m��(�#OI�슀�-��Չ�6��X��j�n3���C��꤃ϫ7�]��)�%�n7���I8ʂ*i?Tˢ-J��[eZ�Nx�5Fs��Lq��o�?��ZX�Amp�NbeY$�1Z6�:���i	ZD�A�?�ꭗ�����wsf��@���`ӛ�*�#@��23�y�]ї��o�4�2������aAs8z�7w���}p�u���H���0�������=�k��T�k���c�O��|m�o�t`��V��-��}� �������:���&t�p�B�AP>�����tz��h #�(�- �������EŠ��?��g�p��~�c������ s9pâ�����i��.�b��d���J��l�NH`Q kb�l(�TƲн����L*�����x���;���ܚѶ��OBH�)SpI��U�tUx�Ҕ��b\%�фE�&E�ɬY�@`���n���D������]6�a�����sb�h�Ƒ�p��g������?Nx�}��A� }%d+���a���u��e���.�������V��i�7�4�vw:%�����S4w���|��P�rpۊ��:��q�rS2���k�<<Z�`�,x��m�?0�18Ȇ��[��"D3�4��
�}N��ɎU��o8�c�pb�C����S0�FifGI_FS�e����⊔�,_C���q�N��^�[:�3^p�`���r8�OJ^:[���&�h�Q��gL-��k�����U�7	�.���E2h��hx�e{{�'�^e(�3A#Q�3������I��7�`:�;��+�>C|F&�u��w��8|K��=�.�����`���OCz��[�~��d�	m*3��^ȷ_�B���=�\Ж#�"�"o�}h�)��4&��m�;�T�����˷�:)�=�_G�������/����M�cW\��3+��w��b
e	�FK#u�M�)�9�k_�9��
P�Y���~~Y5��4��&LQ�+��vxF�4�+ʢ��p��=Bg�e�UL;PwmG0���u��	_�zg% �-P}�>,0��W�����K�=�R����ή*NK��<ڼ�����?��P�=Y��Z��gC�kX��]*I���ù`U�͟ ggg��������!�r'RO��^�
;��hC�7&è��LQD�-L�0.��?��k�$�U:�E}�/��Y/��nͩ�T���y���+�ڦ- �@��Hg����>�z���~�]�>P u:��,~�����ջ_�����gm������~"2�Ѷ�݆=��A��:o��d	����
Ԅx:x��~� H���'BV% ���ߒU�Zy��*M�z���=LII/P��C�������n����8���	aOum���S����g���l���,N
3����R=���M��c:8��,�q���g���������~<v>�p_aq�#�������bu��Z�ܳv���"O�@�u�X����CE�I��Nr���X����2�%Z�������O�\��N�C�꠽��+��Ș��|ְ��F�!��*���fK�W�=>�J&3���m�݉O�T�����8�=��h��~�딻1J �wo9���A3�f��t��'�����w����Q��;�r{�q�'�---@~���̲A3M�P�>wݣ�K�=D"$pj�A{�������^ ��mN���
߳�
0O�?�c�ַ���.��7�,Gf���J���%U��K<�8xk�k���"e��,/�xIx�+h��V@��L�Tf�s5��*�z4toj���J�ފRoވ��ΘNd����:�'�x\� �E�!�)`i@����_��UQF�7�l��� �����~�H�9�F�V]���W�0���k\g�i`;���w�[ZXS-�
u��v�O�c�O��7Ό�����V�K7������뷵��:��#۸Z�����XAT<jݑ~�&�&P܃�-��7ދECg�e������t��7��h�ó�Ī鰫T�I>*ǝiQH >�c���7L���_~ROl�(AsTZ۔�suh|B&�2 ���4k��d��؋��X��xs��*��@���-��>�5Qo˲С/>�2��o 6�Ǡ[�
w.��'O^�`O03�����>�ѭ.5�\�^�}�*��S���6�GRW,��"�}�5�C�`K�d{�Z�t�W����ք(����nƉJY�Eo�,�9~�R@���ɪp���b�ql(o�^a�ߌ��L���u��'�޻��
S��U��]�}� ���9��7m�띕�MrdI�c|l��Z���н���_��FM �|Վha/��r3�XDrUֹ6վ{��Q�eq�� �9LU��#�:4}ы���>w������s�1_?1T�y��W�V�Z�z�h��Жv q���c���ʬ{�Do�����*��zX��Ր�Bj�;=E�UV�a@Kn�4UHh��N�k�.�/���C�LgF`��hD����DC�/��b�#p�J���OZ��?�Lx�1)}�}���U߫���]�u���`���m��C��{3��@;e��v��05�<1��4��o3.&%�Y�!��N|�A=!�=�}��z��w֯�����9�2���wU%@��j��|~�iϿ9j���H�:�/s�`����� �XR�.�[����l�D�� �Y ��SC���9��SAؚP%L�)�hn����C���h�f�է�Y���')�p��^����B���\��W,ڲbnr�$zKJJ^rrQ�4�tל|��K�P����i�O֔�o���Mi�p8��S?��O��?��u�#���R��-4d#��~�-���۰i���,T����gY����$�I��yݓ��;�+p�R�����Xnx�?��
w���iIiNk���sգ�83�yf�g��6^K��2*"�Fbl'�N�����d!��-�7m�_?(��	T�l��:1����}{��y��D]*@Ď�S�m�d$y襒�	#���B�h@h->�y���G:Eg�=���1.es�"�[�������T�Z�԰�w��P�k�_wM��ȣ@�^��j���eM��D��
�+d���JU�0�p������"Ǭ�-$�|�Sl�U�'\P}����FP���Y|�Y�qYx)��͚*ܖ:50}�+)�O�g��0�5A��PZ�}]s�]�>u�i"���4O�@�<�)Y�������t*���l(Iќ���RbՊE���"��"�L"mI�e�����C���Ӻ��:@D����^'i��TIkµ���_-�$ďߖ����v����e�Dr��ݯ�}r�ӰS��?���T�rCjM���J���	��E_���e>�IudrY��{����^�,�Z����o����M�}թ���u]�����6ہxx]m�ۣ/#��t��=�ww��m +����&��+Xq��;�J�gU_ڪîqu��q+���I���G-�6�JԎ$Z�ΞO\ Dm�Td�D���6O/��nHU��e+���[[�D7���x�տ�;uj�-9^<D+�Ke:V�������ĸ���I��o�L���#1������9o7��9���_���!C�R�����.�3�>���_7,V�����M�VAݜ�c0�'���c?v�Wz1J{��m�(%�� �x�u���ؑj���i����mN�Ϧ��V�ҥ��i,BD}�{*C/�h��j$�!��+2�\�P<٥��sL����f��;�o�☿�鈏�_�`�bK���9���w�Od*���eo�}��N�u<���A( m)}[}v�b���Ũ���\��'o�}=e��^�
�w� .S�<���=����x�͆g��8���F�7�:>���;S�5"@k��tJ��������H�뚜4���Jb��>���r�4CD��R����[6�[��'#Gn��'E�>3���L��x��%[*A&c>G&���C�n��t���qg��t����=�i����'5��eKn�Z�H���d{M�p8��������=��T�xw�af�I.˸k�ϫ�߾"���x??(���B�>�'c�2��G1���7,|b#��B���'\֠;��ʻS/��J��2}e�j��(�l�t$�{�� Ó5�H	��~��sǙ\Y���t{G����=�w�՜RXh6ο��,���q;?_��e� 9�)ҕ���	p�Ӭ5����&�&��_�J*���S]x`��le�q�����LHB�K�Y�l��ZU�_���e����Ճ6����>�� ���2��,���Q��ir^�-y]�NW7���`%((��VCY��Ϳ�t��QU<G����&�i��BQHԳ�Jf���:�5E�`;L�tM�/�C�W�$Iox���V)F�����V��l�����d⌓�#�7`F�o	�g¬9QKp��_����a��JT��Awڸ���@,�&u����A������s�mԤ*�V��9�_�wrj�U�[O=�aFzP7��;/	�:���������dX�U�3� }�Fຓ2�.�Y9z���᾵��n"��4�Z'� ��hh�m��}Ι���0p:���mē�2�I�ϾlH�Bh�kj+�ٮ?�2~��"6��َQ���.
�?�4t����q,��r����V.?�9���(�ij�����ACÑ�}c�]���瘧Sj=�j+�R�UA�kc��T�`����@bh�4�X�~�=�t'�u��N��y�-�͋�(y�!�b���M4"Q[CF�u|�������c��vG�h�w�<��c��qIj^k:���KD��w@f�L6�A�������6����-$�퓉�����얆����U�΃]�k7�����Ō�R�"W��<�"��l+�8�C?C^�	i��9�M��f�6�_b������/3q#BVt��hǧ��4�BqN��dӃ��Ov�9�{t�EF�E���}�y.�R%�ʶ�Ҭ���7͊�tו�5E�7~������l�|�ŭ/�<����aP����M�|Ҍ,/g|�o}M�֛%T���c5qʱ�sK�Nӹ�h��ࡎ~n��m�^Ʀ�i��9	�qf_#�x�o��ZZ�0��\_�{X��|3��@���_&�~4��u� *�a��~��!�#��X=��QQ��u왽7��X��ֺO�+����P��������Qs���^�j>{݂��.a0����{}�6�} �ĮC�4ٔM!��rccc�z���I��W)�iYhg�Q\�x|+SUU�P1���ӓ��`8��?$$$<��z+Z����H��JuAX��}x*��|�m'Ȥb�Vʡ����+�٬H/EZ���s��6F`�b�_2�m. r�y�a��L��v4��i��L�e����+W��'l=��o߾5k�+��8�����li���e{��4��2@�Y/g"C��E��7�í�$�Y�J�����ԦUJ������v��\�'�Qs��=P��}�@�g��J�&�)�R�/��������˗/M;��/_�����䟿j��K7X�bŊ�Tf��/U��
��d7������"լ� �k���F��Y���FD��b�ʱTs1x_R��9z���#xQ�֑�qT�1$1b'�9z�<_*yN�κc'�ܕ�����|�dg5��51�BHM�>{��OG�s6����s�	���a�Z�;{�7c�t�e��������8�$�MY&`�|=EqW�����~�����oh05LŜ�������
�,��s~Xx�V�}у��	໑Ɍ�!�Iԓ%w$d�qus���~��=�� %T:��6HiX�'�.o�#�~ͭ�U�qEc��������ں�T�J����j�M{ ~��^����[(��4'�����]���ǍN�/H��(��gȦ�'�;��.��('llk�=�3�W2��~I�!�)eY��[b��>��C��TZ�iE������|�����o*�ne���)�ɦ������A.��P�]}} �s�]�3��|F�l�����|�j��h4�.����k���.�ʹV���B�l�/�qʊ��)]���1�[���ЕaH��妫�4Z�,�_Ƕ�����D�|]�J�rvs�^��Q��)�X�ŋs{�Tj���9��{*��� ��$x���n����l��1~s���A=N�.�xw]��r5����ԨL�w��7��q|�f��)�ԀK,vuCÒ�y�Ǖ;������֤�
�^�z�-�Mq�![�Ls"��*�=��:?���>a�]m�Wr?��� IM1p�A�X �PyWm�ҕ;�f�W^��X}������۶C��ʊW��X^j'�t��q��t�%^QI���.�l�p�p������������J��]^5ң's����S��05q���A}�&�������yte?�CK�$�)��-���<���'�KyxZٴ����v@�oC���QHs���5�!��h����q�H��u�p�e�Mg���2\��;��yxx�r�>��?��s	󾯟n�ݛ
G����������m�X�[d%-����GbD���Qu�v6�\N;� ��a���
+
��t�t×V�p�;0`�^GDb�V�:H��ȣ���]S�����\�p��6�ޱ"�d6Ir?XE/��g�;)��/�����v:���7�"���-�T }�'�$}~���.>�����]<=��Θ��9'�m�%B��b����|?(��~��B,󫱡�����jbv�W�T	��G��5(���Fǥ��;�y�Q���]���Ԯ�{��ج�2� A����J"x��3�u��'ƦD���,�{���uТ�c��cn~�x��Y�i�u􏠧PSiYhT�|Q�?pS�����x��T���?����>c��u@��;�bA���v�,�1G�a$��w� M7G���'���,9�t����	�6s��]��p�c�%3�ԧ�l�7��;m�n�ן�+=q�8S�b�W��U$�W�(`�~S܃}������c�E�`�hd����������pG�t8[i&n�`8��*��U��ɑ�,�;��d�#����K%� ��Q� �%i`���u��gn���'���s��~�����׀e�~���}��D�iNj����)�E��k�͛�:jR.��~>�V�d�Q�$�TtѶU�}�̚��"[̶����9�O8�W����e��{����Hm܊�ʵۥ@r 瘂"��*�F�r������2䇹��a��E'�d�
�f�mQ-G�wƴ;�>2#Ƴ���w\�3��a�bT�3�j3&���7<\�z��\	),��+J�%�����	�RU���s@��3��E|�g�w/W���z�.���)Q��ė%�/��9[ŶA:n[;z��]-蕸8;�p{�}��v�O��W���E- x��-\���!�sl�òD��/.MEz ���ٷo�Ϩ�Ե�s)����#4���a��k���77��� �P�|���q�\���!��A�Pd����Z�٨�?:���bB�<$L�0�C�T�L�.��=t�c����̽���»��膭[̲Ԁb�������a�
���[�m;����
|���k���7���^���W�,ƖE�i۶nM�9�@ >�ROw��rf��Yq���Iv	KmG��n�7�������m�>p	���Y(x���UdA��ߐ���Âi5�E������M7 �<�$��:4�{��~ �G�Z�>>�B�&�ݗ�X��P���4�mͣ`�E�D��h�"f����{o���}�������].&����Y�'��j~�ُ�Q���ywx�J���!7����Nw+�d]�����B&DYEܲY^�kϭ�<UgY�H�+t����9x�.@܆�	�g��o�9y��]#�֜��������K�>����;P�u���"���9d�Z�ӬG:�z���1ZA�B���"�{g;X_so�{�'�~�^��K�_�P}��C��^���2O���EY�Y2p|Vxp_+����\���{s�x�|+;;;N�l�=(O$)�%&�Yn2P���+��T�!��V���bP�-3i�O?���9�!�O��š�T�ࣲ�t�۰m�j���qG(~�Nu���xF����S���P���<g�r��oN�c�m��ץ�(�v�ӌ����M��I9�z�l��4�Fo�TԷe�7�T��Т��x��K�o}}�E�6K
����A�λ)���<����&��m�sm�2(/zy���������G$�R�/�[�0o��4>���$4�^��ө�Rꌭ��U��������3��ܬ��>�l���"I�w%���y_Y8�F���]]�J��RQW�	Y�!��sn郘I���S�B^]ml좹c�U�(W7�g;]�f�UIS�Q���Y�b��Dq7Q��L�{���e�`;�c�^���|�c2�RXe�K<�)���޽{EV?�Al����B�]�ܶغ:�//�\����r�g����v �}pJ��ą�YM�����A>չ�^X_#�)G
J8�L�3m)���Ke�Y�<���TRx��1.>��j��]/^<y(J�������-Z�=��Uk����6B�O�^���kIIH��E�����a�W&0]F��p��!���q^�����)vm�"m��h��e�F=�b2��]�/��c�E��gV��TF)�(>Y�,c��/��S����wL�X:/ύ��|H�"�u[GP@�+�r�6�!�-�ї��Io�ޭ��=%��k�o|3>yiW�E��|Y>������X$d�|v0�h|�#��ǋ%C!i{��P�lK���j�wB� ,}��m�Ԯ��m�w{�� G���m���ٝ{|����n�����k^!z���O�^�`�U]eS�7�$l���Vo�H�`�iS�1EEE��f��������!��ʿ�.��=��b
e��}��z��uSY�,j����tb�TJ�W7^~������*��w�N����8��~�����D�q�qv�@m����=ԁA}#$�mӗ�j7c��S{[(�(����^��E��u�mv�e#���Q��b�Q�,+k�W/!6���Q�Ԛ��1�.�Sh�����F(3x��k�;�QWڭ�M���kM�Z��n>��䍇��a��Z���a������"��7���Y��>��P\Y�v�h�O�����BI��'�����Yl:0��/<����|Z�rS�kݑ@Q=���������~3<����:�K�K�����-�u2�m�.��[*Z����##�u��a��b��@�1�$�gG���3��{��T5��ʹm�����օ0c�
:�A���XH�z��-`���Ww�m�\��R�d�����:G���n �oGh#\M���
�V�,�F���m5����uhm���A�߿Z�OA��}���if_=���c��*��NĲJ���Z�&+��iH���e��e*�;98,]�SہH�8��<E�H]қ��u�]!�ɓ�G�|5�0v]+f��r���~��-��u���u�ZTԝ�ߜ^�ڠD1� yٛ� �5b5��ME��I���nlj� �x��P�����]槒��3��&���aH��E������px�F���t�F��4�PY~�C]�Zr����:m��GU��d��VO�:�\/�$�픚A�G3-�$I��vW$O��5����L�4F�C����É,�	4@��g('n1���%x,D�1w�"�^=�C�.	������q6sW�������nt��s�
�l��dok�"���A�5�,\V��n�w�L�����yEZ���P���1�����ƃ�{xb�v�*NI�SV��������������8&��-M*ij�����ԩ=�B/)'����EA��d�m�|W��Å�Ȓ������}�z@������F��ȷ�Έ�~MuY���#��G�n*IY�r%�Up�cc�8 iF���VĴ�Me�B(**Z����	~����2�#|����,u�
.����i?�F�O���0��u@&����6Ǉ@�P|F���E6���7�{�o?=�3���xT���=�o{1d�l�GF)�w_u&U�P�E*�n�@��/H{sg�_E2��oI�Hh�B }C	�2�ov���3
_�-&[u�R���s.�����ki��7$A�y�'���CaOȾ�˅n[��@��}�m�Z? �1�]=9h��p���O�ff�?��l;.��L�������9�P���L�&�`���ŋ	��Z���U��7];I�k��Y��t��=���r�p��P(�6��=C��,b˦��k8d�=�k�0� �yxxX�Il���Q�A@7K�mI�Jo��=�z��%�Q��Ą�-x5͛�������
t���0�⺁��f�m����?|y�D�Rѱ��;�t�)nz�A8$�6�����h���
�Ào�Y1-T<�Y�e��򾻬���ܫ�K갋9շ����M����ON�T"�ݜ"hA5#/����1��V�bQ�z���<"[q�-�_M���2I�j�S���W �0]7�:}Y�N:�3�0� ��9ற�5�k�]��?�IӃP�^���<�@��b��gZ���ADۂ��ZO ��M��$��h������Z��ۘ���Ρ!������� =��T�uj��&���#4�߬<��7�9���W|���Ŗ]��2��<C���î�ғYL).�X�tم� �2⾕�9Q�,�&��ūV�.�,j�{�2�	k�G����9��:�KD����:��I<�?}6�ś�7o���KdjNL����Q�ݩ�k��\�B&�����kp��t��m��%c�-�V� 5��ccc/��Ի�Dg��0u����8��A�%벗ATH�	E�-�'�l)�.��I�K�y�~�+O��#��8�J8p��A6T�ȳ�V֭�xDA�`A��pg3�.
"N���`N�[ʫVUU%NK<���z�����b>!��z95�ͭ�~��*>9�Zt���]�5��R��H����=����z#��`��
2$,<��,����N���1˻�w��N���Sk��{*\�w�ء��PP eh��ŷo�.d���g���yO8�S�T)Po�O���U- 'c]����ܞ��.uq�ҵ_\8�������g��!�Y�I�p�4�'�ɤ?o����Ҍ!�v��J:�^��<5U_��O/ߎ�塁 �^�܏5Sʍ��&�r]7�;�U	&O4H�9�0*9��<C-w4�z����xP乹��D/�Ή8�5�������B��j�Y2?0!�穦�{-���Ua���r��\o	kO�o��Pf��%�H&)��A����,�⩬�����e��R<���(�<�Et���|�qZ�x9m�r�6$���n��"D.���ݳX��ǟ�?V����O��`����-�U��"�wMk3�����-y�v ��]������ѣ�t�����O�B��q
g��tݐ�2�:�L�b+�����S:�L)W���Q5x)A�FE�1�V�9�?�Va#Y�nA�_!��/�1
<�e���;4t$$xc��e�2֚Ӥ[����hV�_���q|dd䖋����*=E+�n(��Wc�??g�Z *�d�+roMq�3[Q,x������8���)����q
r����9�KJ�ĺ�/=�s��V�kj�0��//�TTR�b)����2�����(\Ԭ��y�]f���c�������"9�W��]dqS5?'��ao�^mS�c~³y�������޺��&;҆ī�I�N���VX�z�UI�	|�T�() Ru��,
N�{ MŮ��9m��z�ut���n�VN,{[qcqU��\�³�d�w���*�-ySE;vhG})�&@5�w?�vʕ��C�Fy�R���^�u���*�v�!O�}�8g�*�#n1������jy՗��ni>�:nQRi��4,:,;��r�d?��z���7�(��k�j�+X�M*��t���� x�}��¢�:28!S��}�ú9 �l!��6��]�@���N��y�dւ�j��N�����a�*�V�b����Uu}�i��GF�j�3=�`�� �E��s�q
w��}�zː� �ibU�����E6q��[  5V���lB\dcS:������+UUQ�+*��a�X ��++�.�ml)O�C��;7�m�K��Y��Aaw_ےy��a���@@���8n�A5�l��֟_�A^��?gfb��aR��t�M1ڙ�	J�G[2>�>�9������;ېr��.����{S���8�d�7rRA6��k׾��f���U �/^��t���Tn!ԭ��Ϧe��_�_t\~h�3d��4���y�l�m����.mA�e��%�)
Ҽ6�?­{�ĕg��b���� �g6��^��s� Xѡ���Ï���Hq���-�Ÿ)NA}����gth��2��]���m�9/W_lqjF?��6�ZK����0F����M�\��k�D�tQ\|�	#�����~k�KL=Ft��n3)�̫&j�_KL� q5��Y[t3l� �՞F�k�����+}3N�)��m0�������I֬���V��76����(,=o8/P�{����(ƙeL*̋b�7V������r�w�5�!j*"��E'�Q�q�v׸���c���_��8��^����r��/�/y����~�cΉ#�_<�bժ�
%�d���[H�����~Z[~�����ܿl)띌Fw�">P.Dr9Q�?���>�-�;�<i��L�����A(a�;�r��`M�Ԏ�ԩ�@�7_��[M��)h�b��N�-䶜V���#�My�
�����Q���|�����bU�ng��9M��}n4�!��E���M(4�)i�[s��W��hѢ��οm-��s啊�"����9�6{�Ϻ�0��}�|z'4�F3��^��^=㘂��Ą��w]�H�x���I�/4|^W-i�gv�x	|�ј��6�����)��l��Y4�
g�R� �9��ǝ!a�������<�) _�����������ܡ���|c��K�J���,[<>K�����U㹭� 'M����I�#f�����z�Ӣ] 8��)�\���h�����m�=N�᱾��i+�Mq��D	u;�Ѿ�\!!!a.կmG!���y��}���Ɩ��ْ;��.��Z��~6��'�:����u�����R�vP���c0����MT��9f��(�
��ʆ-�&Ϲ[�N5�?��<����n{)�"*����eE%BD�\"C�21�iC�d��=T���$�N�,c�-1�h�2��yu�����ߟߟ���u^�y��<�y��I�d��Y�߻a�bt�����M�:�4{^�.��J���9�������Xs�1��� Q�}��V�����0m9|�䱮h��ẶHЂ4���wIv�\���\O�*iL��ӈӾO�]���9�w� 8A]����������G�4��fD��x�i�/��nS��#��2�pK�|��H9i_�G$�U[&k�W;g)Q���t�� җ\;���G���{5��]��S۬��?��~Y���oYX>RI�D�[��x�<F��USx���\ԕ���e�ӰJ/�d�XmC^?*�~G�����s �ЙB�=_��*�JN����n�jL���~�"���p��l~E>Sk��Uҷ�֌d���!u��[j�w�0.�/�+���N��= PMiҮ^ell\���P7��'��i���$x j�\l1�+#Ds�z*1�-��Z�<�y
�M��G� �C����fc�
(#�D=:� $�i���iZzzS?hnį|��?�_��ç��F��e�����d8�F�~Z;��#�7$e���Β�T@�ɛf��zE�$M3�f���a!ϟR�J�6###��~�q#�鑝�N#���?�>OG�/ݿ��E�o;��V���0���U{��Ĩ5%Rr��P�����nn}<'�p���ˡ�fdb"�~��B��G�j�~�&����Ã�J;�0�������5�ۄ�����Iv2R�����Ӫ2��i����,;���
�#�3����j?о��)�yH��M9�����l<h�(�	_��>����o矰�7�E���R�o�D��O�~���0�bo��3��.��ܪ�[L���P*�yu��X /��c��^&���B��_&�GFGW���u�:�|%��6a�XX>�\����|���!FJ��O;:S?)S�$u�@�y&����yc�t�?�� l��u����B������w�jN����N	�|�~J1�s(�;b��9Ǥ��S���c*�R��E��H1�/�����Ϸ�7)��x܃��s�-����r���z��X��S>ף�t��կkM�}����Gt"�5�������O���2���mC[ˁ���\t6��7P��^)�7'���>��= ��ƣq@�����8�H;�a>�ݾ{*�Q8����Ko�k}��z�$]�КĪ�K{ !��-���;�sI�`ėm�>h|�vN����%M/�Z��"�o�=Nn�t7������0iu^��I�������Հ)��P���܌��}Rzv���]�0�.u2�6[=�~�<F���9�֌0$�J�"O�ۯ�o��p��\/
IAB-k�[q��%�B�Ӱ�"+T���p��>�4��7�:;M��[]�ӯ[�_F��cդ���׼MƦgg���*+�,v��o2~�7<�B!ctfRbb!\�n�0�+�U�K��a�n�*cR�l%��5�:WJG�^��B�o?�d��GWD��:���N��jc��	�gX�Pt�&��|��[S�$]�����!�Dk���9|�碲r	�w�T�xow��Iy�a����������>����_r��~�vQ.���|�#O���s��\��
(>�i���)��e]����	��Ke�<���	�:��"��J,�OѨCt<�;p�ضg'�v���y�{�n��.聺�1Vn3�D
n���>����1�^q���_��[ ���8p_`��
����.`���:�6hF���/�-@�0|��o���O��W-���Hڂѫ.g3~��P3�8�A���]�Ky^ywݢ+wK�Iy v��J��Cؗ@�q���ͱd!���Q�����M�WPЦ��*��z�F���l�8kw|���0U��Ð=o�����o9z>��u4����N9�W7��D�Zk�^ZxPf�wF'�DH�e��;�x4F����KӋZ~;�=���N�=d�d˥eu�ʸ��,�p� �@0|-�,�eOo93���^0�A��.Ve�;\&[8qbgH��n�'o�����6Ji���9���v�?��˗RSSs��p;��H��H��d����ͼ��s�y�����Y��	L��&��,qKӁ~Y�!�3N���,�I�
��$�#�>��0�G��N��-�ͣ�U�����RVv�}AV���䴧ha�ӆ������'�~�+}��/�#q����<��.���U�G���ȊS)� �m`�2�Y'˗`0�} \g��P6�����4�$�&��q�h��h�Q���	M��o�5F߾�|������X��վ��N�8I5n:�o��o
�q��*q�ϛ0*��ν4�G7��������mAS�i�}��zr.�]������1�G77Q�QY/!t��;������e$�S(�Ӟ�����d:���N-U�x��[ɶ�1Z7ݍ���~Rơ_敖bB@YE��;9k���?W����:���Y�!F�0���R
��"�'0ᦉ�D��#��ڗyy�4�"�ݷ�Vɉ�I�ɦc1�z�b����ݛF�^��֡��� �R�	���n�C��F쐐(�8����z���ͺkb9���羇䋺���S�!�G������3eɥkQ+W,�t|}�\��j�L�v�\�T�\��y�?ȋ������,z�5���s<��44�LԇXLMJѱ��/@迤���}�ZL. |V����z�����`ʮm�� �C���^T��;�������@	.C,�_'�0�sj�Rp��\��؇b�Cѵ�#�#����f��-���_NLSg=&���C�*l��YtH��Q�8�����df���P���\�YY���~v��V�����W}��=���nnh��}�&�PV	��m����Y�w�N���P4A�w^"�,�kچ}�e�L�7q=G���r����g�h��_�n�0����NCض�+���e_
���^Ot�b��q��\���:#������PP&�Rj�H�8�?pQt��g�p�����K�1gO�3�*����Xt���+<!w!�[�4T>]�$�p��3g�8]�7�%
�#RC$P4�%�?��9������?TؠM���u8ŢS/U/U�Uݔ�����5��ϝ�55կ������`x�Fj�fN�n��+�ؿ���� �n���ﴲ�j.�ptԳ��3
����7p�*'���q;����0]��<(�GA��W��K���%&y4;�W�>��t�S���d&@Z��ؙ{^c8L��j���n)�њ��9�5�)`����ܰ���/�u�t{�2D�)焆$tGJ>q��������V��0p���5TAm����O6����g����s%T]�sa�d�AzW$6.�����������@�5\(^8M�oA���.<r�tJ	݆Beu�Y�g��|��>0s����'����CCe�GՅ���h.�v�NM�����)�Jg�k�p���}]������	��X�$�E��iT���'XgD����-�ɰ���WQQ�{��$b�^�`6b
Lu-�vW�t�DQ���100��*+��#S���.�ą����Rv�Y����T����{�T����Յ]EI�3Â�t-�
���Yl��q��0`S�ԩ��^�vb0�V^=��:*#������S[m+�E3>J�7��qc5�XhR|I��g���,�r����F�s�lv�����l5���B������xH%�g��xN��B��R��]���D��'��i�o�Ҧ5�|���Gqn���' � P�z$Y�_�qqqy�j��_���P�M�/=���sGr��b��<o7��Y�Ԅl�����TF���\#�D~��I���_�"*�ՖbƓ�w��M����C��~�ʀ��]iM��;:�*+�C���d�s�ٽ�?ȶ�U�Y]����?n�s:
��������6쑌��+A����"s����B�p�:�(6�ݬ��nz<�(�Q��U,�9__N��ZO�$�j�A����5P�f!���,��N6g��K{֬��n�UX p凞���2x����"�����c��C�;�f}����(��xV^d��O� �_����<��k-��"X�DN%�����(_��@�O��*0��,�t�DW^��y���I=,�l�-��}y{tt����fJ�B
�T�@������
�!Eg�5N�/���Q�Ҷ�8cۑ$׿��a8�W���1��I/�՞&7*�����W��	*N�k�#�ȵ�"h��k��k��D��N ǃ
�1��[���Տ$MgQ(��
U\�S$�.�����e�����o�D��?Q�m���^Tg�e��b�LT__d�kv��VA*��8�׸�ĝ���y
�ыa��?]�C�"�qM�%x�S�Z!PSRR�8?�憃�Y9�c���{��&�1�7���j�g�W�3m|�[P��ȉ#1R-ǒ��Q픦�&�����~c�Y����LizP�"�^YUtV��]^3�^b�M3�!�����#��+�;��e���
㒨�����9�O���l�bN�GG��/��lL��P����a#���j�վ�FN�m�rֽ)�i@���y�5�Jg�/:���e;y�JM�I�##~���_�L�4�H�#��`{��'���#<\fr�6�����Bu��	�w֑�}c{.]w�jW\���>z{�
�~III=��U}�N(�$j
���\�����jc����
Y��`G�+�6ZTɝ�Wl}�>9�� DJ�����M�*Vք̓l3����Ti��G����N��9��as��̛��Α��
����P��F7��ћ��t�����\z1 {�����1�,j��H���|�����:V�0��r��$���ϟ� ���~�>(�"����9��싷�vm�����2�~Or���$�S�z)I����%.M��e��Ӄ�{G,:�-� �1��ռ]��%�R�G+�a�hN�c6�w�8+��CW�Ķ��e#k��53�J;�[183kcgU3=�Y��ڭ}�g׉m_��:��a|�ڴPp�iq|�^�6�z�OT:899891�X����k8�u�_[/���#+��ι�ɺF�i�m��$�\��jY�=�������3Ƭ���}�RE\������j_���<����ˆ�3=�Ś�Ì�I*I�|�lu\�������ۉG���נ�P�V�M�Pg~;s#��۷ĩ�����E߃J�%+)���]�|���]�d������������{C��1.���-'-�Lu۾i�E�|���J47�失��m)�7(�zO:}��|f�l�K��u�xPp�I>vQp�,�c^0�m�g�,�> P=���C�\�-��m�k-ʦ��tE�W�q�F4vV66MN_=�;�	����`�dƛ*Wx�A��*)J�%��m+eXd!ͣ��n�N�� i���I�"]�����[�d��]iBUhO~��QV�7�1����O��}����'��H�,�-��g�R��$�NO�q��T;�]�j��#{F'�h��6�S�tE�S���@ݧX�+��FĽR���J J�s��0֦����F��u޺n���pKx��xJҏX�F%�l�%�P&�Qx��ۧP��U�{Y��{��4
5j$RH�l��ϋ�D��<���"bp"���4	?�oo��#���_�s��������8������_Cp���7
ʇ�����V/���i���U>L�!�}]�|�-�I�Pb��[���~z�3(�H�٠������h��F��@���r�n|X9�Y�Q��&}������I���$��Y��ol��0�����ni���'�h<I�-Kc�}��[kW�?#`eG$,��9��7r{�=��p�~Ǐ�忾�r���>��j��9��R�^�j	���������4iII����-�iԱH�BZQ�ً��O�t�-d&�+ʌh�����_Hg��w(�ZdS%Z~kΫ���&�bqk� -�T|���b!ؙ�]�[�sff�R�!�l�r��]Z���S*����G{��N��Ǣ�׉-�X�...����T-"����������1�������k�I��Sݖ����pp�,��-H�XF"'�lXô �N����h'�K��Q�ߍ�?~�����	w�7n�MY�`��<	XR��j�!w1F0��r�*�-[���Z�Q��&
G���3�]c��$�>��FvC�����v��f"��zi�����A��L4N�av.#�|�~���Ç�x��~�
kHѽ�4"�k*Ll�%c0�̑J��/_�(�`��CC�٤Ǌ�{2�����~���3sW��$�D+*8�!`�F�Y�+j}���Ƈ	6F=�����{���\���<��"������}^�o�_ً�3�M�Swm����<A����R��ꪪ2� �p�	y�]���1}#Gxѻ����T��OM	m���{_;�ɤ[!(�-u����7֨�����Hzƥ;��|d\�y�}�X�f���Ѧ$��R>�[� !��Y�Q\�	��a���M��Nx�M�H�4g�7����n�ϰ�a��G'xmp.����)��jKIF��uD���ԓI֓���7�� 8m$���J�KI1�����J��LoRB�I����@..?����PK���q**����&�q�b�VJ����k�.5XvG9gX��Ɩ����
��l��E���@�M��h�����v�(�o z�mV3��Xof]LLL����F�!�g����r&�5�*���� �lWfgW��M}�ǻ��FC�4}Ksww��	<���
�>s����q ��6~A�@�L�X��v��cI��O?�:�������9y�ǰ��q=w|�S�Ǧ�6�B� �y�>.8�tM�̥'�A|���D���|�yG7�e�J��&����ϷK�G�1G]�/�(�F�cU�s�b�nL�������6>�X�o���'#�)�H�mi)��Wl(����6z����;-yJ@Q������G-�R��NS�1�-�g��~�ڥ��O��FIf���{V,�����J��/%��zۥG�ۮ���{����Çw�7�F^�~�֍p�9�3�F�D@z�RO��������~��X�C����ѣcۻ
�'F�2��Uk1�d�/�^Eʖ�C��3zF]wr��c��5������Vj*����`[����7��FEe�@>|Q'��,�����Tk\n��ƽb1@֩i���#��q)�{���_����@�
��5�|�HE����ݜRO����,�x�G���`�$�ʘ7F�3�R���^�ü��֪�����$#�-]Wt�A�)+ C5�^�-&ֆLD*����@�+P՛q�n�w����D����~W94d[�ڢjMu��n86Y���^�]�?]�΄��o=�0�}V�����̷WԐ#}�)yV����s�!b�������"y�-�3v�}�M�D}��V意y���YGDOP>�L��4m�6�R����������+�H�5�Pz�t�J1�W;�ܹ3��\[��S�,q=����V��j�١���=$ z�����I�%���W�����<'�_�Q�V�g��C��,!u.�۾���Z�D+�3��9c\���� ����@,����y/-�����i���ǐp{ݿթ� �١��z"��_Vtmi����h*�����? �r�!Ah�t1 ���%��!������C��HFd #Y����(w�|��|�C1P�[��&U��qJ�SnD�QV���&;'�Qж���-u����(�^NT����|�|�M�|���5,�EΥo��T�J&�m���Zܱ
?��6yZ"ɇ3�6YF���E����K߄���4��B�]�R��<�S�EB�5��lͶi;p�smDR[}���*ɑwʜF��.bv�ʕP��'IY�r�K=zTW��,��r�*���i>���!�Dj��H���i�O܉�g�T�&7ɋ����~`���ihh��5��^�ύ;!�����]����B'���6����,�y��>>��e|��Ύ�������� `x����?C/~��fPntS���>7��zD��4��a��Pǖ(Cڂuq��
�̅ޱS��RpP�9�rqf.}k��o5'���u��:&&\r���0�q�['C��Z9��֕1.��m��u�a�@ �?xy5�m��Qe\�Ɏ��N�)l��0h����PxIq��o��5$����!+Ev�]�'�_�M%�www;1�H/��UWlO�Y�ϩ�H1ғ@]l��e9\�<l^9���ع	��_a\�E|��n=���١?q7��`��/Fv��`іmmKyy꡸�ۈ&W��Z�=��Ӧ��P�&�Cgg�E���B��δs�?���0ZEZj���97"H-Ο�5��ok�5:�>���?�5��mX�H,�����
���8��B�ﰺ�y��xIEE�]�i��ȹl%�3��K# �0�e�"�bݰκ���n�Q;���3� �U�$�S�N=7ю�waΜ��Y�� ����v�曤WB����ݞ��YRT����A+�����?C���E+��z��.��T�PO������3o�jf1�@ڜg�,H���<!��L;���?��|b58����~�R�bȈ[`:�-^�O/��s`����|Y���B%��7=���a*7�T��v�'M���Pm����X�E΂ȁ�H|@w�ŪTl�72c���#/�vb~~MY�ͪ�jk?a�(V2H������.h,�8��d��?�ȋ5xN�t�W���^������'��OϺ2���L��A~yW�'đ}�>~��3��z����d�71��Z\���c����-�C������3.[V���J9��q��!�`���uc�(�]Q��WPṷSD3*h��eڜf<���jq��
E�R����ӑ�~�����Ր��
����v��g˝���Q~ ��u}��lKqZ�Al���xE���-C!ok_���_��
A@5��?���s	n��!F�[h�y�W���`P>,B��L/����9V�6 �s�^��ζ�3�|�f��`d�B�==�[\����IR�~�]�"��g�i��k�
6dZ���~�Pwh�8�&\��>ho�ˉ�(�!���{P3�'�d�D7v��h��F�$7(�������rnvf��@~��UM���ʐvT"�'�t����i����a��w�����C��2�k������ @�~��*r��5���U(���ar���%�]����,����&�$�_Z �u��`�gQ�Z��Ģeϙ�wt���e�m䗒�p��_�Ȫ�t�sqv��>����s�]���L )S �V�(}jɅ���2�]%<-����if�S��l^c4�s-A;��46D�F�F5�����3A=%�V��b 0>:!Ё�_2߿;�h~��=�1���.W1g�׮|~���Bގt�Q��[�~�N��7�fG��LorJ����<y��Z�V�H#y��&��p8�9S��F�X�q�-~�4���Y;������;�	5v&�g��*���N�������e��'}Wo�h)��x8|�:��ğ�jqO$�N;_���1�CU:����Q$|�����9�� ��=T�¨�J������6F-��4na�Xr�U����lSP5(��.�!8��A���k�~�G%%Gć�Cn��?��mh��ͭJ�A� �2H�c��ƶ�����^^xY��t�׾Z�?��?�����0@��C�ߚHZ�5l +��Bw2����()��<�#g?vc���犔�k����|?�s��+���'ι�}I%	���u�ۺd�?��!�ʣs7�9�R|Y*�-�ٱ79�.FEë�7������xL^���KQ%�.k
s��+f��vD�[$���q�Ug��΄}�4��j�[�b�G�D���5�����`-����T���/͂�w��[e-�E��yg,�N���w�4�� i}[���j+��w� �2���.r��PN��"�"Q��gs��痾\���8��i�IzK~9�c���W��?�"�9�g���#O�55�=���=����-����Ha �$ :��G�]2���?� c2Kю����L:me��@���$v�^�yuռԟݭ
Il���F�:�f^��As����]��㪐�f9/'�WV��"�w<k��lB5	8�}g��%��i[cg�y���b�#=��B@���Y���8�ؕ�O^޽.��>����)Qp���ha2s��ݾ�����!�/��C���Q�m@��&7��Z0���0�#�&m!�?�H:�)�!�^z2�0�e�����ש4�������7�[?�^o��}�¿�K�'�M�y�q�}ci�OY�v���
���x:(P� ��e�G>�
TL2/�%��Ӿ��E$߿�����[��L��Cf��	�,{s�����o�,ܺ�v�P�
��h�}��@!AY��v+����ȑs,UoT����S����c�`���ՒԴ�����@������閿@JZ���]����ӄi��8����ȫ�݁��Yd<�oRZ�J��_�>��G	�q�\@���n�e2��̿�?+'�*j��j�d���$�C�7ڮ�/���u�K[��<����5u,�/_>�و����i�F>�+#]g	�)(ճ?L�O�Z~5A��HA��k�����؎�t���k"3p�h���ge��\��ƹFY|"l����{�79pF��	��?��,�gh6�ni@M��Xi�l��[gju;(��P��Y��eh��܋ �q�"S����a�1Pb��w{Xy�),X�$��.9�ׇ�R\~"����e$��w��3X�yA�K"NU��y�Y
�x��3YU�a�j�*g��xN5��Ν��~�Hb#��"ը��r�"�L/sW��"���~C���?��i��Ov{�鼇�E�	������P{0;3s[�S��u�z-��n.x��j��A���?�V[���Px�^��"��(O�c��EC���
K�����ș�_�% �V� ���}����xrncދ����������|Y��i���i/΍U4f ��@�����UPfN«.b��!��9EC*�f�\I��Dc\���Wuy�q�%B=G��H+�T��V~4*8s	�ѽ=
`��*NN?��K;H��
�<[1�:���h��?q�[~�	Q�dsC�9�Q�'kZ��f.h�T�L�۫�rx�ĺ��D��h�X�5��r�Z&����ļ�`�ҧ��SV�hTH�iI�o�i��;6���]��<���5ʁ
|���J����
��LOYY�ųgkRT�Gcg�M?֤�RN�$*R��n�K>i�(��[ � ���ת��q��{s.�8&�����W;=�U�L<#��#��S�a*P���n�8H5#�B��~�U�7�f��O6.J��,4x��=z��8֔��������vY-��/��Aa���V5��X7o{�겆KY99;�����{W��]u���^縇�g���vR�'V��={�A�m�Ҙ�4����V}��䟕��FZ HO�iw1��C1�QU�k�`Xt�xz��.ϝ&� ���K����������3c�6� �&�*��� }��J���_۽�4p�/ ���&p�����n�@�M�$3nKH<�ӧ��#��c��"����m<��0x*E���Z��ɋ60׿
�������|����c
��Tw>�	ʴ�nn��Z�I^�p#�������4���s�<)lrSC��W d���%��G�h���I�5I��P ϻ ���|=�����o��U�[z�P���҄����A)12@��zג�ݥ�ڳ.��U�#2w��/|��(Ԩ��k����3�������FA1����+�s��𲡡3�F�������8�Hv�^�[���h���;����w��$FH�����ZC#Z�(��:0ڔS�$�ӽ���k�����:��k�;��hlf��u�[T"�j�W�|=���4ע��5K��E����e5;ׯ`��#R��IK���gdB\����d����4��?�&�~��n��Yj	O�I`.��(}4ZM�m�ȼv�?�4�䭉	��.U���Dty&}����;=��V��ju2�A;<�UGc-wh��, {���/R�����+@�~�ǡ�|46�����*�I� DR�T��p�x=B��P��i3�����:�D���~�w�"�Pjg�ͼ㴇����i]�T��&���i��36Z������b�[Zı���hS�='a���1����۬CL��̑�eOU���������ꯍ��ݘ�J�E��A� t����=`oqc�%�:��0/�WZ�Ѻ�E�x���|��]���$��Ny|��RbZ���G0��hB�Ma	��q�̈́4�C-�Wb��%�n�?��r�ͻe���K: 8��O%7K(@_RAAbW4�6�d:\��P���s�,���S)s�%���of�ؾ��=>3&�����E���rl��;a��Y������E��ӟaS�-PC�m�!.6�4�i~z�@�ha��@����ᴜ�+�c,\�P��(�e��ۧ�������
�� �϶�j��N��Ǡk��'���+��V�^��6�=�e϶�V���^V�G��Y���C
~	˦�#\r���S���tQI��u�*��0���	�3�aA��3g���e�����Qg<M#BV���p�k֔���3jl *�.D��Ed����!k�gl"��<|3_�t��^ڑҔ\w��>g�.���V�n�X������#M���{o�"LG=ۂoI��?�@�̛ر�rX3����t@	(o׺EXb_�Uc���B#���[��;�GO���d̵$�_c�R*���(�<�=��U�}��HO�$��Eh���ڤ�E�N��0�#e���ot��}�~����y�W�I_����t��'�+|)�w�7%I.nd#^~�@:�N�����I���֥�ڕ�_l.����V���	�d;/+���r�����*u���-��?���)��j�"�i���'&��&�����޳y+rX�����D��
������<�<��A��3��-��:ǪUl%�S���¬x���g�1�hB�t�7tD��m������dن�M�kW�!�|�><&�Zoq;̆M�����m=���"�~|�4$�;�n��>uk��jn	x!��?e"ǣ��v���W3Ot[�&�<�npQ9,G�?�aGe��ȣ�kYD��z�a�{�����\���I���H�7!w����fy��U�|�������H�k���঑���ԡ�}��x�55�4w��j�AvTk;���pE�#-2���Uc��D�C'%~�����J"�we��dز��-x�t���{B*��e-��CQbn�IjdDOW17b�R�}W�WU݅���h�oGL}����Np|�EGl:��ձ�G�O[:g̶��œK�}V^��@ |l�[� ���`���U���4ՙ���[��ˡ$��F�%P�u(�9;;g�n<����=���ʄl�̾}�۴��w�ލ�_�W���d�1�E~b|�H�MbUډ�M�O����j})�t~L�`���_�$�FU����h����T3}����Q�0�z���������7���R��D��y��@�_�#�k������]��װM�zL[ ��Sz0�SK S嫙���n�}z��l�~�z��}�`���C5~k��z�HXU�Ƶ����֦O ���9*Z��x���U>��}�������U������()��b*�Ǩ���>�U������Z�)~�5'rX!����@����i�O��/P�������T��<e1�0O�(2���� �"B�t������$YK�?+�;��=�DH�bz�^��@E���<;<1��x&V��o l��NM��[��UW�\92=�EE��7��T� Ϧ�j�7Q9���ׯ_�r�����."��t�g�+p�?�C��\�qhi��Z�l)�-s)�"�x�%��rQ�x3������Q89���I�s=DCs�]O���V�˟'޽�m�UT��D������W�=̧�m]t�D�i�"B�5T����T�C���OD��O�v���K�WU�:�"���PJ4f����tdS�3/���?ga��q �/Z/�d�&�g�� !݇�T��+U�{�Ծ�*��7վ�� N���d�>g���7o�
�]�Lv/S�sq�9@P"���*�[4c(��D�'�j�N�"6j]Cug4hu�����@������nl�ڗ������#^V#,a�Bn�h˺��m�aT6�9���_�fQ��c��u�|���P姳�g$G�N�$cI�ӵR���
Ʃ�w}��-5��C�f^&�O�5K�jO�����S�Eօ]w�n�<g�#�;"�NШ�J1k����.	4/�A�X�:š��,�z� ������F.��Tx��F���]��:�"��rQ� �V)���G�_��Rm�J�����Q}�.D��qu4�O-Cmc��E��xMCɪ?���,�#~�������\Y���ׁ���G��d��7�=L���]�-�I���0A'V�}SP��6�\�z�\�&
g�r����_�9�����t��<���M`���v���s�%��Dʷ'g�̞�V��a�im�n�2̀��_8�X?��y�`l�p�NsIwy�jp+�E x0���t���e�
x�G����K{H-&�#yF^���������K�>2�RN�w�K:N�ŋ4v�~y~���Y�����A�y��+;�Rɷ��}��0@�cF���g�B��^�37j�f�
�ь3m߻kfK�C�VV��3���Ӵa6i� Gz+���_FWN�?%9>k�aB�� �� &��r�#��ќd����D-����V�L���c�a��R_NL�j�EDD�W Ȩ}���s�'�غ{���Ǩ�b;>�f��G�dZr&�$�������m��vҶ��;lj��p�X3iJ�}%){2�
�0�μq�'xm|W^��O�!��6���v�O�gg3B��3H���aaj+�}Fk�n�/�b��j��iA\���= ۾�QLt��m&xW��ѣ���
��h}q�gf�YX����YQ�D>�S ��]I�u�\d�/��*�h�-�r���a�TƟG�-��T��V4�Z~Ja��#���9��cdr0Y��i�тf0��:9i�.y|�M�F��f�[L~`�*0������f��0�[�v�� O� \�Ab���v4���`�Ǿ~Y�Q3s$έ�		gN�!7h����Zow���P���	i����HԽ����'O'>h�Y��4r)h${���c=ۛ�k����CW����>{ b�M��@_���QD�su���kW�s�(Y
��$iDSȄt(���ٙa�v�Nև�<�Yd���������ҀJ�K5î��:��#G$?���R�Y&
m��)�Ǒ�U�gZ{���C���X7������ ޤ?疕h�#PK�q�D_xo$��~h(/��F����54*�	�sĠ�/��uA�JjHЬ��8��$�~�K�)féP���o�d�_x<:��AO�u�iWO�5>�;�V��yy�Ojz�@?[��;�6���@�-	��j[�)�]��	W�O#(���h��M�o ŵvs��`�/���\ 
933<k�BkC�tlk58�E�˪6*8z�[��������T	i�sl�r_C$�j{F]���w�[ڱ�"�����Q���� _;��i\x��JD�ד,>��"���ץh7ۊ�Fr*^%����xI�4;r�x�Yb����v=��W��y�ٱٙ��jPo��ͩ��i䚹��V}[Z*>���A�p/��vM�yeZ����m'~��S�gQz9{O믌q!�EO����`t#���N��Q��N�� �uK������~�=pQ/��K��G�Y*_M�Of��L�|�fL{Q�/��U���r�moE0nx!�A�Ͷ�8CtY�,��Х��%��X��Q\�q�#ׯ��;��6�������ZD��I����b�U�얕�d����(��L;���$$�ep�2��9i�˱[@st��Ң=I'��NE`{��y�g�5k�:�2m֝�˙�e��������H��'�:��ɖ�*I�N�cuaEF\''�q̿x�@�J�9��&�"R�IHj�iCxP�o��A�
��=~�a��\,��%�z�^�0���.�r�M�!IT5���nM�75R	��� �0pb�u�F��������`
u�� �G�tf$d���v�̲����#m�l�-����6�޸�P-$��h��1ɘx�u�[��;���4��?����D˟���D�Ъ�����)����m�y z�"����@�*�2�����ck��wuߺ.�H��>���{�g�L=zt�LY>@�jͷ�|G���F��6y��:��g%Zf�~���Y�[m~���RV�׌!=I��΃�ԯX��?Q��Cj�|)-��1c��|	Py2a
��:��T�CA��	|~o�{5��%����r#:.�����T��L�:��+��=�rIp��I�4���9�_9����NVw���=��@LLoeH�|���g>��/��r<AK�V����c\�1��W��Y�ޘ&�H�&��V�N�m��/�0�w#�	@�\F��ڢ�@?�xL.���>��f���s��H.ܺ��fu����\g��ҵ�,ZH���Y|u�tȔAQ�da����#, ��H­`ϥTmJ?�E��~��d�A��#����7�I��"�$h����B����>��[�J�T\Y��Gs��f��l�3�m��*Y��F���VW��ղ�L�m����߅ΗӍ����E<l��ࡀ�i�Y���}���nKck@�m�5���䆻7ڮ��VFZz{qq��$j�~���ϴ$r��~x#�D��mV�4������$`��MO2FBk�߲!�Yx��Lc�a���Xߘ��v[Gj�%�gH�8<��e�q�?y�7��ƛ�_a��/zrv]���e��[�&����ӟl���M��C��S$����*{�Q3]��sS
���S��x��U=N򞹣3�L(��ݾp�=���l�;�'�T��Lo���}�+������=����wF��� 7�������Ƭ��a�3z��)fɝ}���>�� �'Cg�H�P�$E�~|���s���'.��IǾ`�\*����6�|lI�1Y�N�&�H�^��3(�̧��E�%�I_�����L���nD����W��t�ϓ�����~yY�M�@W?H���������q|�D{�߮�����p*,�ȅ��1���}�m��|tF�P��ɱ�ضA�qn����Y�����@A�\�b�kו�P��jՠc��ԩx�=rGc͈������Z�j�nt��}ɓ���{�����PkyktIGr��iw���!=t#��ro"{��hK�T�M��Z��Z�r���K����!&��k���Y�j�B'
����o�����ㄆ���3Z���C>DK�:y�}}}��[:ˀf^ºǷ�ܩM����ؤ���ˤ�H�K�YՔ6���I�U�:���J49��H4ZAJHb|�6XF���:�F��N9�<�蠟�_�2'�ͦO�9ty�wo��K��l�@t���Q��P�����-V��3�x!�c��� U�S��N�1K���b��[f�R����G���m�Y�����Gጿ2ܚHP?o��J;w:�%I���-�R�N�Ҟ?_e&,<<�p��0�p��0h��X�ܯ��uK}�l9�A��|acm����W������*���J������s�V.�0�.�����ڱ^w]Xy�ڹh��`�2��p�;
���QR�Ղ�~�M�m�:�²��u��/�����Lz>3�LA�J��������Bᝮ�[&>pz� ��{����^��0	�]��$:9��ūM����*�߄����l�hnTB�Gj��W��[Go��KXB�,�_h��|>�4����/���P������bN�݀��(���������3������
W�ߔ�~�Pg�ͨ8;Q{�ť������ɩ?������AF� ��A�x)�o�uLL���<��[�7<���|�#_J�`x��W��.~��q��?�Ƙr_�a���=��6�9Ռ�_݋��>W�`K��5�P��@�%h��:7��X �9�~"�d�-��ƪM��-�s>۩W]ֹu�,<=;�f����S���y:3����9cI|Rpl����V�B�][ ��T�K�h$w�ɮ�+��(�9�#q���NS��ʘ��xu����A�ml#}�z���ɪ:j�M����ipn�i��{��9dm�8�0u�z�������wPv�����?\m>/Ճί*N*���⫝�w!`ѫ��w.���*�CHq��K�ō�AK���̝�Q��KJ@_,Dg�����M"����DH*��?��@x@��6��$��MY�*�rޤ�\��aWW�I������]��x�~�;np�G�^�W�3�O�cC�PFmR�S����'��ҿ~%���
�����/��w9����� k����m�^XEPQ��,�0�d��l!�̰i�UT��f�%�d��"2#�	�%#a���@�O?�����ӧO��}�{�k�{�}3���"߿4�nڛ�ڼ6B��՛=�e�����氶m���*��ϕ�F�Xǜ�Ҟ���5�65������Q���hyi��������������AD�U�ي�3�.�"�n��tGȈo?�����S�N>k�P���lo8j�'l�e����s��W?d{Oᖑäķ<�k>-�C����^��W_���?��n�G��8؝��M1�+��A�w���.������� Y�k�=rl�>w$��1�`�i�T\};ޠ�����c�m�H�$+O� =.)됭���P1	�J�d=�A~�]�j���z��6<wg�W�t���s9n}{��R���z�{���f��iq�9�U�!jd���=pU%��_�zzX��+?�O����n0��
�k����5?M��f2hG:g����QCT��UO5Sy+D�t�Lg�Iu�qX���X��sE���[^���	�b�������/��F��{;��Y�Y�+�pu�2�q�I���z�­����	T���RP%�>W�&Oy�� j�☀XJ������
�^�+���2\cC**4��ʸ71Eme��������ު��w����v>��2+R3K��yo�sh�>�(��>%��J�e۷J��Q2+71ڂ���e������"�wD���i��7�n:�t#q!j�����/ǁ*���/�����Y�����'&=�]=vYJ\kN�¡���"k^��%&�B<��U@ȅ��Ax��;�:��v*��\���~=)5]]��ƶr�PI���Ԃʂ *�ѹ��)��$P^�4�8�V�p�BS�9���A(>{T�4PE������Dg�9.���%�a��A��5r��F�/�Eh��l��։r��W<O�m͵Az�կ?o*�N�<l{��KI0�@%(�]l�uBK0I�tv�t7 ��i���2�>Ƶ%󆡩3#.��ds�1�kL.�R59)����K���	��UO��n�S������I�A"['R)#$u�n���{���2���
g�������y�m}1H#ʄ��\j{����C8dȔ��4�;M�ߙtN�yj(�]1���mn 5��c���*��Ƕh�Z�O���S FQ�%7�I]����#���#a�. g�%~��r�ϓ�CQis�ߢ���M��J��,>s[#e\������h��F$Y76O�l���T#:裕��.���RO��I��Ѿ�-9�Xx��3<*�S�_�i帏���f8�	����ϕ�Ɏ㳾���-�Q	
�B;7�X!�Ikxj�C!�t���S�L��R*�[C��w��'?��v2�Z}G�3��ZKJ�熊�o�G������f�g�288��-1�8�t��]]��C���c���se"u�`H����T�?��Z��_���8j�הi!�j6G��������\�tA]V.��:��̳hVj��ԱP.>����TZ&�*T��?��+((���>f�ľ�b�K�=�N���^��WS�����/B�?02ֻn�
y�!tuA*�<�V�#���G��ݎ(�R'\| �#�4������[�j"��r�)���ڑ�+W�k�	�����z��8����`�l5����Pǂ�mv]]"��un�V�Zv15�7�\A���ua_�r�ښ�2t�5m+:ٳf����~-@��
��OYE�X��%����<��^Ӑ���H���o�^�iB�HG���Z�s���E�5�!2�$�l���HL����&&`��(�1�ݫ?��CU�ta����չ�rB�����v^Ea���$_�ż�Ǒ�+����(�c���3ʱẾ�w�Y�y�{s��<���Mjz8d�Q�	X9{ ϓ�J�v<�.mp���c���|x���~বS�جl\ `�q�I��^$�˕�;Kcw8�E+z��/t�U,X�`k����4��+��>�7�#�f"�2\�qj#�}x�S�2���&���"n�cmo��_��/��$�^�"��WR���}�UY�Xn�c2PQ�'t��J_�.\�+�����c�	��2�Q�$@Z��˴}G���W��7{�7$9�負�`c�ٛ�2���� ���ٗ��S�t�N5�X��|d^���w��@N���?pL�m��u�����8������W�����r���OQ֑mۘ��%�D�;�6FՔ��GξLB]�����_o��#~[��%����kWWSc�N`U�(��~͚͓��#��U��=$N�ޚ��t�ϴ&B�I~e�ʒW!=�ʮ(��
^,���]}3�0�m�~�;��� Q��+��H�ڋO�	�~�SD�aU�樂�WY�P�#�u�r�G�f���F������^�ۺ���9�fЭ�.�ȷ��B��J�СCH��'�3�>�O���^>�o�ɳ�l8����]F���|+��������=3H��|yЩ���^��A�d�
عv߉��6��(�ׄM�nL�� ��(H|�.�_,����.��Y�����}�S�e�oG�e�]%w�nn�}cp�����X*9����n�_����Ss�Hӡ B��Eo&�]�YВm�#�a��?PqY��E�C=�������ns�~(�Yh��@wbW�\Y9�9�:�Y�}�Oo���T�,���(�G���mgg�B�;`��!-���:j�2���+��QGo�ȯ������(��☗�O��ixQ����p�Ko��Ԍ"M�H�ӂ�<1�^���(a�=�[)�G�0^�	Ȃ��ti�>� �u,��LV�kJ� ����ak���{?ݯ�m��7mfdj���S]ʄꄍ-�g��i�0;B�E,���y����t�f�]���l�����/T��?S�W����5��� �E��777W�h�s�tN�g�<���G������4>5f��Ѱ�H�y�t���1L�C�$�=�$b��#�cvHl)�k8�n��U�-���cOͺ�U�.�ƭ%~�8A��;�716ִ�I�Qq�xk{;.�vC�7�LQ����?5����و�S���mXSVv�;�56"�q�I��|�>��J�;�P4��hL/��-��@lH���q[p�����Tf5Z��SA�����],�0u|q~���.�����Zۦ�� �mD�c9*��("XjqN->�w-�����k������W��:����L׷V���=�-�� ?�(�����.z":����F'A�����cee��	�f3!�8�g^1�l��̫2��Ϗ�Hk�W
B��ȥg«J�7r1@��7���󟉋Rpפ���Y��k�xD�.׼�>u*��/���1Ѱ�Y�+]��o�J�G��s�/���uz��3�u���r���!���ǵ�k��K{��r���mP�;�(�]ASo������t�5A�96}�,#y(Y"�V�7�:�0#�����AM��H�x�����<�o�lC{}^��Z�ͲZZZ.H�����:�P��vN�=���H�I��D�
�qx�`�x:;~?���W4�[~` ���}aA=ڱ�]>E���g��������4��~�Rq�t�C�yp�a��?�Oç��V���f>w�g�7u]�Z�~z��ȏ��P<���{���͠)�D�$rŲ�-Sӳ����[�2j�5ǥ�z/zD�'��h/��񔿆���+�M�}[�����!?]��(��F����/^�|�c�?���1��ǃ�� �ܽ�8غ���	)���W��-,���N��hE�\�X���t{j�ۻ��O�/,#�gR�,fr��Σ��4s�1¯ԋ�OS/�*'�ρ~�R	0����Y��@���`~j�O��3�L��@�;���T����S?�@��_����CK|>���B���ǒK���^���Ӧ��N<��ZOK�n\HW�-JJ�R&���v���`�t�>}���OF�n�x�G��m"��\�F7���mY�f�?��M�iҙ��YW����ۗ�������mw)��{��H�2��x���]�&=�5�ѣ��B;7�ƫ�,����uɱ�/�d%pa)��?��	����.�g�����UJ�$
�b��xVZZ:"&�9���qz�%��/_Δ]�M!��}�騜\25�i�lk���������Gz�D*��x��Z)��%T�X��6���>�c].����I�RH�GBh��7��G	c���4�l$�h�w�M=���M֥�7o���	Yo�4w����d__��@r,���d�kd��bWi�Z��(;�X�*�Վa0��ޚ�Z���!h�Bӳ��&ߛ�d���W�0���iR8���v����-v�(N9r1��g/U�.�f�����B��S�M�J�+��{�+��>P�OA
y^��+�M1�V{Wh�Z��۹qh�7�$z)�}qUbd���¾�xNS�x������,��ﱶ����?��M�.�����w�=o����I$�ْ�"/��III��56a�O��г�a�-xrB�.jK�,��)o�0���^#0N��U;�	�jr���{v�-(�ZױrJ$��t�����E��իǟ7�E�,n�u�M�)��i���x�	m#Qr���aͼ��˳�g��s���RL%R�	��k�C�G2�
km}zi&h�9� ��\1?�ڼ�nƪ���'�0M��h�a�'o���x�p�MN����+L]��,����������j��ˢ�5� ��tb���w��m/?�tt�ґ���'Z���B�/Lt�'��a�R��腻���d����/���0�ai  QRr򆹧������VVo�|Q��;��=�>�QKr 4��[��W͊G]L�$87�`/���>�
���[�˧�W��,��Ez��S�&���)�Py2T5�n8D����S,ehnj�ȃ����=O/%�O�o*����[�:�u� ��د��Co� �F���־��I�4����(��^w�#:T����!�yy��^O��s��\�H$��ǭ����ohh�[R��Y�h���8:f�~��k�ȉu3�66�`�ubB�'�/�e��;]x��L��"Ж���W_�
�Rh��W�:�A�\��d#�w[����v�8�D��L�U�RLR������́�U��b�l[s��͛��qU�w�
O���=�H�0-�j(�y�*y�����߯�]�7�Of	���P�Cw�dLV^ŷ[G����ȉ�O���6N��4y�1Q�N�+�r���ɱ�.�'��sCs5N�ݯS�o`--U��&�R��C�Q�����?Fc�g����v�V�Ap�լD�+��a�e��r����Q�����PI�u�E��SO���ݛ���Ѷ�GꙠ�n�=����rI�SFEEe��t��pojk����6��G)/�����,�wN!�i�i�-1��D�p��>����Y��0[�����m��L2�!��c�� �5*::�Ɍ}��?���Ȣդ�j�63��Oڢw޻�*�8KY��h�G�@�����Ez�bM�<��C!_@�7"Mu���5���ݻ;h&uutt*Î�����u�����V�y;5�a�<�H���^j�s����vz�䋂�n	t<��j&bN��a����3���'��F�����>wԍY�}8�L&�I����puk�K���i,N�N��)��Y?�5/m���7gZ4�V��+����Y��Љq*�����Z�K	�-�?��N�[�������Yf��R��ƴ���o��}$ā�[�=�����ѝ009k����Q�=��?	Z�K�S�^����t��6#{_ U��+w�(��XK��h���&�珶����Ex9�QϺ���C=\���Vt#?����C"�!��C�<�8.�s�ojN��&q��K.��F�D87��n��;�YZ�L��%yW����Y�n��h��0O�t[Z�st߰cs```�K�}	���S������
�uww�$^e5�?I-cYZ�B�ײ�"ZP?�zyG��t�]�"}̪���#bZ�|sZ�W�3����Ix�]�<N�qh׀�[����S��FFu���%,���D�\�:1m��Q���6�]{��(���$d��gj&^9���Z�j�A��a��e`�ls��߫;�����	,�,:K�ok�m��x:~�_��8�\�����DoSz�#R�aQ�!���n�3�i��=�vց�w��mV������B��U��A��H�'gw�!��t:���b͌��u�VH�0O�l�au��&�_K��d$$p�Ѕ���z���e�۷oG(��A��O�Z�*�աa69�M�Sxш����A#%���{49��&��p	��`E��*���������7�/A��C�?q�r��sr�)^�5�m��گ��=��W&e���D|��!J��ݮ�ql�>��3�B�0����<����h������ĄG����!H{���I��t(�Hx]�m��"">�	|~���[ʸId��E�GG?|��Qά�lG�B���F�Kan�e���M�g� ;�}��",��$z$���>N��3L�c\�����ܼT���gų}�s��tT��!F�mx�"1??�%�Si��׿u���C/�@��یfL�>�Sh$���8�H���0R�y)�3$W��.�� ����z�����ͺO5�g�T\�8����������.��6��~rn�!]"##�a�݇��;�>EK��:�^=�d	��\��#H�>
�ޥ��w6;��79G��z�'ƕ�"��h�Y�*��쎸��֚3��iB�T�烵�~i~�9)'?��E��F�#�#k~ġY/�Eg�%&�6����ΙgH${��֬=�T���6��0xԙ?z�^�B���3�XSAG�����{Td]wp�&Qp7���k�ж��zM:��^zw��fE98�1�wn�����_p�ȁT�E�`�3XC�� =;�j�N�M�>�1:K3a�m]]]��v��*gn���1Q���xs����@jNnn���k�ڂ�C���"4؂P���7|v��d�Fg\�HU�_��}	��u�U��q�@-�VF�<����tꉸ?�j=�-���s*܌n���56^H��@Fpz��9^=(7/�f`����{׀Q�����e�t0�x�b�m����hg��;�@�V���M4{��n� �j��ex�^ɡ�8>e
z�ς�)��0���Fe��y�[FTh!,~QW�f�[��m�逥���h(��׍5�nV�oVc�?444��.�$�
��ȼ�⚓��z+�/aZ����(+����m�WWW�:�KҠ�ޘ�;�@{v�-T��H�!�*�p�I���xo�l�:;�(aml��H�i�E���S�?��'YE	s܃�zЏw����,p�+z��׬Kö?1k�1 �8T�������?�.�mq��Ilm�y�}S��Ŵ�Dx�L
�f�:o��ă��c��P���!�u�����4	z�����%m��r.���d�MM��Ə�8}���
.��u襡ѫa��+�67�^t��hrOOO��~hk�`NO���u�P�z]|�iH�3�孥��/G�ـL.
�v'��ϱ������,�+�!�@���>VO�m��w�_|b�J9b�
!z$%K�M�C'��F
[�RU�Om���f`m������G����/�E��:��=F���Ԕ����5��7��,m�xil�50�UUU�������ߝ�v����5��h�@���!�t��)u����0!]�mN~DZ��Li�D�%�M� ��pl߶�;���"�;P����@�W$[���� �����λ*�׬�M����w������ݻw�cwl,=�W��;�^�&�l������ �[�"�/���3�¨������u�F��L����!H��L�Բn��n����mAX5������j�t�kNkr\�%s��\����F��\�mMssEM��D29�&g`B��U69����$�H.��j	��W����]�T�9">����w����݉�*���ޅ��n))#�����e+�&5:���uxT���wvu��Du�b�c�SRD�
��>n�&�CLOG���P3����ϋ��)���ʻ����B��3c��h��X����.a	#�FQ܎�T|����K�9���5D60~�YV���h1b;G�ߌ�@-�ȵ���l�R+{6~*'�A���9�X ׶��70�yx|a�+@X���?~��� �e���X��^�#F�zeW�4?��n�K%��}�HAUr��j�_N��3[�/���h��rUj��YR�@4�7ǁ-.)�z0�a7H�J>�݁M�{�C���Ϝ₼�O�,���)�#;98�ZՔ7�����(kf��y�됋�a`$��� g�GFG�'tJ�?�� ����WI琍�ZN��0��>兘{�����a�=��txk�÷uv�̷��Ō\����Q����Vo�œI��̓i�,��:Vw�����B�
EE<�B��
D�|��H�Քݫq�ŏ��;9���ZIA@�_�� '����<�������iI^�(��g�]
b�$.���M�&s��aگ��'%4qn�P���okk����[��S��=70R���#��f�7�M��J���WAF�0Lm��pI��QMTDD6�&Ӳ���5��_�y���Gڢ�MU��5���㛍_�=F~{�&)��� B��MM}�f�%�c;�KJK3��7>>>x����Њ�2L����r��	?�IޕW��*t��� 9�3��s�E������M����N���@�G[z����\$��΋�κ��������͸�-�:�Y���u/����u쏊� =���°�ō��Kb���ܛ�������l�v
�C����.��N��`�ag����TQ�b��f߽y�����k2i������J�C����?����OD��{7}g"*$�[�^U�/bE1��r&a@d|�/�+��ۤ�������V�0�/���r����^����oߞ<p��Ҵn֥P� 2u��^�z�ݚ�R�.�����Ě
*�a����@n�Oo֥ ���p6�<�}|�c�c6����L��E�bk=��듔��xm#[��?��W5>֊�;��R>�� 6�fxE4��E��H���v�.�j��@�����h���e��{�]
�U�4o�����q ���3|���khu)��n��C����<�db(Me��4����H�fyg����&�AOnFo�'�_$M��_�xdy1挳
цY�r��<߹�mj�3��Dkjjr��.R�������Qy�<�?�f��
�����R4��Ljϒ��_�/0�a��3~�w.AO����� E0P��76����n��)�PZ�,�g���1�,{68U�X��q���+]�W�����e��k��2Ll�)�]U�l��G9�R��pY��4[�=���v��?P.U}T�r}VC�-��,�}ҒAG�� 	�f,�����gǔ7��f�����k�~������tp��C��Ǔsd>�@�1�Yݟ�Ÿ�����(=�'�����&,3@P��K��N�p����U�.h\s�� �u��*��k�����%Ju�D�4�I�<q�:���	�60.���BhD�w�D<̹a��JL�^�pH�V{��-K<d���GnA��Ả"��;���G�tQ�������q������s�8�|XCS	ʶ���m�A�^��PE��1ī q���(�H(����xג�j��W�M���S�][ŝ>��۾�iW��\��A�oV��#�!w!T�\��q ����^��ޡ��^1�9��
_��=Q/%�x}����X;��)#Lٕ��K��Nw���?�#�J*���~�|�0�<�9���{��>{#��<|
R��q�Y����|�kzǦ6�_�� )Dc�#������I���_�7�?�(�-G7���?#���MWƱF``av�����F� �����\ɺvLz�=��*#�V*��r��i�	<i#��i��`T}��]=�5M��}4ePhj���~2��(;c3�F0�2ӱ?��A�Bti�dH������tDJԺ�$�"���诜j�a�`���La���,��Cx��r�kI��M%��i����	���B'��l�+`�����8C�����s|y*��IL���G>����0����x�ܹF4ӖZ�3��i��rQ)��b�u�$���Joٕ_vaM&�\P�΋��nׯ_V���BH���k�m-�O�\�a�+)�@J�ă��ۖ-��\3ҵ5�Jb����J-a��H�%��S���Ң+{�?��L���L� ����u�(Ȳ����ؾ̨R�
�1U�TVc�n�ԗ����������{�%�F��T%�cB��&���_|,T�Fu&c~U��ʨ���Kɢ�����mT���$Y=&T\5Hm|���@`�Z�y=��|�����`�C��:k�$�	h糃�ӄ.�f��X�ب�;u2HlE	>(�,,�l�[4���>O{j���tSh���7�eb�ߌ�͍o[#g ���<Py��s9������kL3��w ������c��q�q�)]*����}����I2L��P�P��jѡ�WZ6�Fsb;�)��;~�L|�U��ۦ�9g� ڕ<c�Q�3�q5�4�\�t�S�/ݲ^iyd�Ǒ���޴+��`qYfVs��<|�@Nl-����`�<!H�_�n�)c�J��#�4�K^4����)�v�*����k��M��֚n6�μ����II:�J�+Ј�4B��P��..W����RӤ?���m����Uk�� IڴO�Z�'Y��Q@.����@�0:Y#�����l�S���ݯ<�
2'g{AK�X�|f*��RXRkjy�:��C�d[�o����_�{R�W��Q9ӱ��}�O?K޿}�(ao�I���Q�F��xz�YOW��ڏ��DV�� <l���j�7���>o(pb���݆A��zyAn�dy�=�������������	��~��7��q��������djƃ�SB�4G�.;]��C���9���������׹k�������Z�֧��\����3j-�R�̾���!`?�� ��Ԭ�փ�g���#��KY�%d�^�sм�^&��غK�l��t�VZ��G�ciY;;����[�?I�`\1�򺎇$ëpD�w**����`��!Ю��:Q�����?,%fJ�-Ƿ�k��[�$ja�(i[���p�؝x�g�(�#!z�7�l:�m������Rߘ�?����"���5OmD{a�Q��<r��
�����
��H�FM�SE��z�J$��3����,�܀v<���d��D�4�.�B���b�ĉ��VR��������^�1N��y*:��մ�4Hc��Y)� ��)TX��������SGCS�Ј���3�1p�ҹ)�ݝь�t5H"��-hJOt9]��˷�鄛�<1��NMz��S���o��Ib����ϏXǱ٘��`)�TF��3� ����1�Bʹ#јŞ��N�M3̬a��W��͡}4R��+~��$�m��Rh�$K9�o��8���":jQ����՛�ֆ�q��ic�	m�vu�F�#���$�� �p�t�tt��)��Dʺ����Z�����
���������J#o��z�	��W�Q@��=77�g��O;SX�u��;s���"�/L$�L�sѢ˶J�j��&��0OJ����:��0��[��;�y��{�ʔ���@��p���$	�KJ=���ݾ��[��y�H5�$	'C;	V1� ;&�ҿ;�,�Q]��%c�X��؈��^z1�Ϣ#��j�pn�`)U�̜v.�&}����<���J�W\+ExZms90����i��	`����Aփ��t~�`g��L|�E�4����Bdd����d��%|-���������vrÆ0誎���j���V��B�����O�:�c䈺m:t�}T��x��I��&����SG�rN�y�C�G��2�nI��wT�B!�T��^<���7zi����1:ȩ��򔯑t�p�/�A*�R�I�&&��^�/��v�(���C�n?����>j�ϥC�:� ��5@Rݘ[�a�8�}1Oڢ	�jY�F�X������!������\�K���L������_f��zN�.i-����̼ �Ǚbʙ�h�s�F
k����ˇ��J��}$��L���@"\�U�>1�Q�up�I7�{�u�}��\�M·w3w��ןh%~&���<0Q���c'�Ν#�� 
;#�@\3����ÍT�I�#:���þ�7<$�N�U\���|~$����w��2���}x��ݹ��}�{ɳ}���V�1JA[����jQ�@��C�c8 ZH񘫔�j��l�1n���J�oo��2s�� �|q%N@�͜�	�-!��N-���j-�yd� ��V��- ��k�u�ʶ��+����Q@j��W��O��i�y�R2a���Ul��`��#����6*��siO���������H�<��J�*!���~����v��fS؃� �|��_ĩ%b�vl�ǰEﭸ�Z)~�!�g>�D�J�`��� E�p������ds9�7rb����̘y�s��h�s�0Xu�U�vtA[-�w���:m�k�L�S�0�()+b���؜~ä��	�N���z��r:�n�O��ÛJ���7�g����;�s��ՍD�](*����'K����(
��0�y��U9�b�$Ā�&`�@Q>w�.
`��C�~����i1~�=�"�I3�S!�2<2bRZ��yyFcaF˳��!DeWx�F��<�$�5幑���Ⱥd�4�l��j����Tm��ԢG��W�����;>��h�]HLL�����kum�7�l����$���5G�ZoTd�J���3�U�ǒ�	��ml�6������+(<�ė��������~�1�L噃�V��6����Es/�`r�����jk	u�U�O�*��r֮7|V�/z%zx�;&��!D�����,O����rh�!['��#$�#9��KpĶ|*��E8N%�}�N�p���3GZѱl/�?@�C�r��+�A]z;��kN�B����o���B�zE�
廅5o�sms�揪ᳬZ�/�r[W;^����-o��`�ZuW}�~5/>��jFM�Q�p��S��1����R�h���'_��Mٱ�[��VQt�c	��kǦP�,8�Ef~�C{�UN��F�C,�y��g$q{=H�d��n6��f�b	��u�����E�61�V�ވr�ZL�ёG�+MT������~�A����C4v�	ʰ�c��{�t��6]-�aa�8)9Y�P_c�DN"������.{JKK�}�R3�p�����倀ιi0&�66�ء�c-��#P�$'L�Z��3y������^(�w|uL5=.�tH�%�Qf�t�0�Ęy������z+w#U��q���k�Z�\���b_ޏ���@�Y�鏠�#j��`i�׍�������TBe��{�m�<�<L_�m
돲=R+��KLݻjU��
+"k���?�����t�'0�ٚ��̕Rw���hק���~9��y�ߩ�(x�jOŌ�R�Fs0)ŝ�ͩ���f��/PA��.�4��;P3��`���v����8m"����&�����]1ݶ��Z
	U��n�u	88���M��ѳ�$��H��	HT�~s�lIv�oUAGG���KR��S� �r=��S��d���Vl�H�� 7��1�Y�lkp���	��5}�J�)�ó3��^�.�ğ/��V9��FY���B�a0��@�ݳ\¸�!��׹��6������Og�4�X�P���E^����ի
F{a�D?%ȗ�d��{��}��$Z��!�
ؐ3�n�]����;�C���4ix��ٍw\�� �k� �>�Zi����1 �e��-�8���@����+r٧9�Bzu\]h���Ō�����q��̶�o��H6��\�_��;%��	�m��O��Q�E����V����n��Q잛+�?4��`>B�6�*�X��_��&�"w�W@IYYY5e��26_��� ��..�_C�<�`����Y5w����co�G�m�G��M���-�J̐1�3N/]3���
�;�%3�+��o�07m"j�76K�#�a�;�	/Vӧ/I�0��������]�lm��}�6�0G��.��wBU�dP������}�X|)Ϸ��0+J��3R>>>�j��1�H&�+�������-�9U��7P����Gw�)����{�x`4ǻi�.m����	���O�=�]�چ��8`��c�T{y�2�����Lue��!	���O��.6����DE97�Š�e^7:2R_Q9��ԽVSa���ĉ�S���@�<�~�Æ�� M[04F��hk�b��h&�Yρa���K�M�4�H���҅^�C��V��er�~n�-G�O�����m--{f�u��2��
�ύ���_]u�9T/ZUo=�n��J��!���r��������#�T"G�p���+J�^�GQ�O�H6LMD�.�U%��j�:�����zVK��WS�Y<E���q�,l�ހ��j����+4@ߗ?��Η��i�H=��7�m˅�B��Fּ�$VT9�Ԉ��E=��W ڃ�O��iz6���Y:R�Z�ڃ��[���i�,�^�h��sp �(U����_����قu�J2=��w�_��eI[v�K4!�-�^6<�Z�'��\�������%K"�{��Ka���cu�?.�u���Ů��n{NSe��z6ُ�i/K,)aT��&�F�M	`@�YZ�A�|�̟�K��p��K-<YJ������P��9R�P.��\��5f,�[c�|�T$g�D�
�u,��3<Y>�]�Z}�1vm����@(��]m�V|���^��5���Z�/֗+��A]g�Lf
��&�ԍMM'�W+r��cY�X�A���&&&1�ڻ81L�R�2��(����i-��sѤG��ho6Ȯ�7dW��}�˪PVJ�v�-����r.�� �ҰB�R�$��L��B;7�1[�
N�U�u��폵��n˗�d�*��vڕ]��fX�A �	���X9�|�eI�D�Hv�˲Y��ve���U�'؝��Q��T��&0%%zk3zѸ��,:ޕ��A��΢g���WM�ʀ�N(D7Q��Ҩ����9$Lg�Oz�=�-�Y�}���i��&M����b	"U�[��/b[��D��19P�@->�LÑh�Q������m�~eߙ����=����[N�=�h���S��V��������;�ߘ?(H|�II���ˮ=G�cF�k���,W~�J�:4� �h��B�9��g0��k,ޝo�M+�F�^���Rw����ˆU1�.���DJ�K��[�v�zWkw`��K�F��%�W��� R��O�������������<�<B�/�RJjSS�\��w�:��^M�?��Ρx��L�ֵ���)�$�� �17?��h�͛W��bg�o���VR�r
��mo�_U�l;�b\�VWn�q��ܪ��\Y_�kbR\1��#���A��/���juL��[��m_ծ�)��~L�H/�&'ejj*�l����K� (%ED7�}6u��k?���c>&�}�
tvl��g���O�%+��`�?��F ���wgHy��S��.��8�qQ�R	��C��W�����QS��8�^� ��^7;���A���u��=��%o�����4�g�@Q�Q`r	�������+Y3�Aw�`=���3(���:��W�rC��=�CQ�r�g� uuu��Ґ���@�R$��L��cݴ�Bd|#��W����h�<n$��k�մ>���ӍCSY"D�i���Rո��#-��?�jI�7�f"v�4�l���0[[Gs~O�-��۰�-X�B��epp��:�k�ѭ��ʙh� ��!��@bvGU0��s�4��d�D�Y���eW��wo���r #=1�]n��������6�
�NR����>���IH7�A���kG�!8'6�8;��M�=�_�n�y�T���h(����7������sf���U��_|Յ��n� ���k^#�u�x�[��	� l��8�4�3GhtC�� �d���m��$«%K>�[�TH�����*Ԉ��w���Q;��ZI�uE]�}W[�%Nv����e�n����}��Z�o��FB���&�ǔ��z)��ࣼhR$?���"^e�k%<c����s)�]��WFu�����d��p,eޏS�#X�P���D�FP8�ي�z��czـ���٦�\;��֤��\"�����^Rd�*�E&�G�;��-\�H;���C����A&Zu�	�3�r��'���H���/��>nMt�ީc3�8"�� T3�|N����>���+-��̧�s�Ks����}r���H|��O��|u}�����D ���q�\"��u��P��\��J���F�uxI�+)�T{j�	M���eߘ a�ħv&_k�U�����R���.ک2�H�y�
����
F��¢��!<O����`<�;|t���o,�U��bk���@�($�=(y�_����ID2sȝ2������2�kkNq��w���x�u|ka|V��ߴ�.
�O�
V��`��Fgkl��޽�<�?�J�d3i�C��yt$凱��u���T09H���4�N+���:/���?"����p�����>�V\���@�������ؿ��B����Ht,w&��C��Ӱ�"D�Oh�\�6d#/�N3�4�+�'���$1Cj��OYӝC �N�R�}�N��g�R3K �V��Y�:u�u}^�4�8�K�XB�)�b/�U���3vn�:�'��<�$�����!v�Z�KNW�-_u���hgQ"����.�F���1ÀP ��x�>�rߍ���x��ۙ�8]�7��n%�.�#f�N��u�F�ѱ��oO"z瑞.�k��>h��K��מ���b�˯�(�Co��[﹪H_�S��G�3&�H��8:�����.��{�:P^F���ba�6l@�8>>�ao:��joXʢ;�ω������ԋ�����z�i�,c��:��G"k�� ����U�b}mot�d�7���(�c�&"!���<�z��qĈ��/��索�A��޵)�.�~~fn�999RE�?�P��fU�.���>���9|�:v��r�4�YSss�\�4���hc�*tnd��9{��D
tQ����/�P���os�ꃵQ����ڸ�}ҋ���_�g�-l� ̂�K����{Q����o��T�+�[���,�\��\��w/��"+�#P68����~s��x��,u�����4�^Dc*s-�b.��'ˣ*��c���@�u~�*�]���c��J&�6Z��܏�����L��w�l&����u�tg�D�K�����bݓ����i ��3��m>�uI��pI��]��#ll�Ңϱ}��<�=<-�g�^y������%�������!!S�f(Bj�FFꋆ���Yk�����zl���LL\�$�U�u�N����\W��n������$Y�׮����C��������6z���'�����i���dsP��,% #1�p)����C�4���h��J����Đߦ
$֣�ߕ���#��p$�s/ڕ�޿��c���?J@ߨ��A��D�k><H��nm"����F�C���K��Awn����qE�T���n��)?�aq�Q)���ח����5@��cJ-���������V�͖��^N)�������U��J��eH���#�.��Hm�w0���
�H�-��'�F6FP����=�ϓ��𢏌�x�h���;�����|ϧ;I�q��,���P����=�үn�@����]��>k�X� ��>	)	l��,۸��$N�.��Ѥ�^�O���Z��x,���p|���B����Q�	m����B����2{�������'<|��pH�+��S�L���i�7��ơ�׬KՀ����8??��N*O╬��ʺ���Zѐ��f�=�܍k`��Mdv|��j�E
����H��!BmQ@@oW�BSCE^9o$���vM����.M�BbQ��a, �����6@UË���Au���A%tL_}�Ԃǜ�Bzk��.��w�q��~�ZY=��j`������}���.�x5�k�񨦴�jF��E�X�	�Qޠ#�g�G@Ф0����I��N)���������/�͡���+	����QK��3}�:�:��
c���Sb�� ��'+U��TE�.�
�3[�_K�ЦFa��φ�����oJ��J�������.\.����ɚ'c̗x�0_�[�V#+]+5���o��/�+s��@ЕD��e��	����x���k@�8�#A��&��Ě~�<��G�QQɔ,]�c�]��W{��ٕ�L���d�0���1m��ů�&mˮ��� �_���_S��J�+P��t����Ԃ��ߚ��3�WJ�[?3����Վ))������<�T�6<�y&j*��O��-��'UX,�T_��;�2��p��m�H�dnaa�K�0�5"1Q3���p|���c9c�9_M��#������������ ��j������Ă MAA�ZA�D\Ddi�i�%H�  �E\qi���t�^P�RX�9ς1y��{�����X�s��{�{fΜ��X���E��k�'^�`�')$���c���a]��xG��@��'W������ƿ���-&|Mf_������v�I��G�����D�M� ��E��Q��������|͟��9�R�"�����]��e�q�Ͻ,O�~3Ū����(<���4tu�}MP������R�|��X�1�����.S�����x���Țz�]���� >\=pBc��R�tt�%Q?�;���~m
�T�eH�w��&0%����h��ۉ�F�ԣd��p��{�et(����׌"Ȉ�Qj�����Y��樫�nt�{Њj�DШ0��WMt�~f(�@&����JMq��A"w�T(岹��<(��閺��@k�7q�gi�;99=����E�;e�Z �c�<�N�k��.�ymmт�#߶/��
��!�����I�����֕��MNN�q���>�~���.�s��&*j��u+�@rO����`B֎4�����%P9~�`9_&|�O ��5?�! �dcm}U������]�l�����!�&G��	_C��_�Ūcw�� P$�s�7�e�Ne:r@yUz�v�~T}�a�g77# 2�sc�yl��ᅅ~kkk���5�Xخ$��m\z�mNk��$%-����Ȩ(=��1.����Y�� nF�{4���a,�� ��I����[���� ��^�xI����u�_Z�MΫҰ���Qş޽��q��^��|�3[�ηX�|���Xm�����K�	Rd�Z�������	���-���~�J��#�&mâ���E�Ip[�:2�E�������M3��-ȱ_������.��m���6?�KIII贝��l�nrh���Ocl*.iOY������#�,rDj����D�Fݹ<�~�A�|���GCOSN��Q��gzO�����?�$G����C�'����:0~>����`�%FR�u]�!�%#@\�J����.x겫��c	��{R%
f6>�\IZ¯l��^*7�B�d:�V�@ôDx8�ב5�>ǒ��{�K�ѹ���&������;���6n���-��x����T���M��Ol�;��T�N��r�(i���C�ш�2Q��B�$F8�F׼ij��9���R�j�nQ˲％��H�hTX��|�]4&�ekG1r��nmaq��dv��%��]
�m��l�;�eR	�y&���+aUm2gV�h���"Q���z����~�nO�I��t�"R����Q2ލd���q�ٞwu�Xqq�(�S����b�ڮN.f��a:�yrH�f�x�2�_'D1iQ�B�&?.,,�:cd�,yc���N��\{ �8!��n����<�zR��]�\��qLp����G���MkTNj'�j���ެa��(L���h�Zr�>�p�P�����&ܮ�m@�Е�{�z��RM����ϒ�3�?��.�P�;�Tw�.��}\�&�H/V3���0-�-@L���d��dg$$$x�����������qF�V�V�.<:19%e��6U�.f�����c�����R��OG����0��vn�ֲ�M������Ot|�]~�@�Zb�]Bj���O����^�Nĩ���zIu�J�{���զ=H _y`��=gt3m���Bxe�j�'���������a�S���(#�kX�,19
7�G�b$$$�<p���7��b�z�1�n�P�+Tqȅ疢���`J�����h�m�C�Ŕk�@����tR6�>�^>�1��8�;�`G��a-N�B,��eV��,@"i�̤fb #�SəlNWכI-��ϟ5�.�w9�7lڴIQ1�W&�/:�ܓB,]���g9l=�����W^k�,Y�1;��9��nTAAA� �����hp�X�srWtY�����h����/ s�qt�i"�D0J�E��^��I-��g���dO����N###ަ�N��}�K]�TCA۲���j���og��ReAt��hHܻ���¼|�n��@��&YW;���@����ܫM��@� ��[TE3*�d!��
���������{)�M0ݰ���Σɒ�H�Æ�(H=1.999M,3&:�`aa�5LV��J~�L`��]'�g�Ʒ�zCV���Y%t'�f�+�um3�����-�<����G�uD_n�Cg�7�\RfFia�V~���1���֛ockI(��2R0[��%�X�g{����e,�o�?RrI%6ۮv�k�ֶ��;���q�������iW���ķ�:��y,���x��rUH��,�Vxϭ������o]�f�^u0�7�A7OQ�R�x7��;D9^�3ח�y�D>�j f~:f���Q���O��R*��h3!��qW%�����͉��S�e�(��j(�@�W�p5�6�?zc�3�pЈ��v"^^:F���(���#�*ε�(O����d/�m�D_���H�a���n=D��J��.����<wJh
��mV�c����u�Xr'c����A}ck����o��hߓ�S�pӬ���mU1W���<(`���#�Q��4 ~�n�o,��B<��yQifD��0��(Y���>��e�wj���"��-�����yt[+++���N8dG����v�����.�h�ʨ4x#ο5��Uv%%���^���I_Gr�Q�}����)��,��I璼�-j�����9F111�v��L'尾x�����H̫C˚��T�
�����7��
�*M�q��bI����S0N���U0�4������;Qυ�u󅴞k�^Ҿ�"ɻƓEwAGz>0^V;�i���z����4��{c�v��z`a�f�.��h(^Qg�3��Z�L
�����(��;��7m�~b����Y����b��������&��<��c:��S�� �Y�]��>������t�˸^^
�!4Bg~�n>A�|i�/�z�}�H��ިpǎI<�����`�Q��{DcHHH`)�W1�zz�S+T�fdd�ۯ��@�:�Y��͔Zk{oU�1֥!��L��K�ԡ��_�Q��[놌C��"l3����Uй�R��t(3Co+ơ]+�_����21Zm�R����p���;~�׹�ޚ�����6̍~��+����O!c�-	))���j&w��9γ�b��e.��u:V@D��1Gm�"J��e8'0Z�ͯÏBz��F�>�%�AL������.΁?SC��,��s�^s�h���#��{6�2�P�,���3�vjQ�E]>���PMd.��e�MP����i���N#<>�;ڬ*`w���u��燵C|R\�!�u�E"�_<���EKx � ńX	��B�"U�)?t�<$���i����4�UTRr�I���e w��1W4�vv6���q��>����:��-N��	š��Ɋ�K�����M�j��GX
��/Td\���:�-� 4�סR�'�*m�6��;�����IeS��6��n��|(�=r"�f��T :ɒ?��7��܂k�L2[f�:����]]'"""�[֜52z��.ݾUCu{���U�N��Y/@h�@h��u2N�pɻ�U�A�75�)�4���K�%5E���<�ejj�pu:���~��1�u����W��(�z6ӶI��U�D���T��?�LP�"*���A�nn2��A?1��I���6�r�9��uz%���ϗu�<� $U�M�.�jЍ�y>Ti�1��P������I���.�3��(&�,�&�Z 5����i�A7X�.�B�/a�����IT2�=��w����!׉��槦v�7 �ۿ�ؙ+|��'��`'(��z0p�o�-Zk� ��+y�)�v�Y*�`_�u�!S1JLw�Y��k����yO�x��1󳽨|���v>��u���P8�ri��(� �Z�:���%��F1J>�SQQ!Q�LSyՁ�σ�X>z����e����j��6�� EÜ̹ �JW!� ^{�S�V�<4����1 =����NBDB3W/$\�}��"�O��I�����_6�׶O��F|Qe�E�T����$�e�w���H�V(�g��^�$&[?ZD���6�#��Q���Qg%����o����(s���(&`u�M�Z�v���������BXF	Pg�؈)�:�w"N�N�2Ag��y�<�;yy�~_�em��5}*��Kx�К�A���Ϭ�"�_����M�@��:�ju`�A�)jA%��Pp)x�M�ncR!�v�E�ݚ�p��Cx�p-�q�B�#����� х+|fQ�J`�222/<�e���1�(����@��|��]z�Mb��
e�P_�bf:[p�P�r-�a"5��X��%��Tx���E�@�(�ۜ����5�\�u���]g-i������~ff{};��.���Z��	/D;���? �B�nmd熩*߽^��������^�8Q4���+�;���)Gد���o��q��n�ޔ��#]f���67��1,lK��bo�v���edf�,"�����~�/��Mjݪ�J�C��˷H������4+8��+�wm�jW���z��y�5n�֫��u��ϻHNN��%[X����g�N;��56Gmy	K����'&L4�f��w����,`@sC�s�O����ܞ��޾�9�����zE�Y"/�����dbFܬT�[,�}�B�'�e��aE(Q��75eH�5�6�K�q s>�������� �W���%�s6kx��"b��Z[G2��FVρ=�T\\��ܬ�X���TG 9�eyv�+!���[�}�_��;L�vsu��c�%�-�W>�§4���+���{閳�p�Guuu���%#�p�6�t��淟��!:���u�^�(�����kB�Ov;H���~�k#�7!��Q�^���l�甪��^g�Kn%�:�E{܎"�����k[�v���?���sHLLq�=�k�t(XyXO��ۭw�.��ASB��W��{��<�PCa����oF���-zi��_~����#�O�I$���;/w�*�ц���"�/��ݗqa�L I�}UB฽a�u��/w/�T<�5��>�do�.��R�W"����d=`��@��M=�X�y1�s�x�e���[/n�g޻���sG����/��2Dj3�^72b^���������&�[���/��r�������+_"�_��@��mm��W/�##k����R��)��/ ��[X�+L6�ӳ���d4:{�����մ��| �Q���'of�ŉGai(Tcl3J�z�����Jug�y����^):�[SV~��Q��Y��iwR�CRn��v��j�ú$.X��C�
1�egg����%U��t�śp��)�M1d|ʗ0�^GxS�'�6?�N��If��$���p0NoB�匒��KH��ݿ���~?o�Ɋ>�E`��r��5���#����$Wi�/����
�WOT���b'Ebۣ���"��ٙ33q�ק1���)��O�b���/ڑt����h�_ѓ������'5�F��wQX�e���8��zxgt���J֬��=�Wc�<�o[� �^SS��2ttv��I�K֯��4i߉���,A��R���
%-[��Q���{���Em'%7/n�C�h֋]�D�;|%�X��˫}���Z)(]��
Nx���g�<3qO�*�vZU�6��*fڬ��@�2��Z9�Z���R|"!4w��?�S�	(���XNzk��@�
�tE�ȒK%$:�1.��w�jT�w�[R�",2%��N�m��]�GT�@�F�n餖�Q�5�����hb�ò����ƮW�Y>��]��,s6�3�ai�'RW���x0l�K��- �8C�ń�'�ꉆ.��SRR"`UZO��
�����9�c	�,_9�D+���kP_���M���hF9X���L��� �/�y_u����-�MG
ރ��~c.�z��O�	�7�R"���R�"��}��H+q4���,��
|#�;Yks\g��>P����z�5�#)#W��� {q3��(�
���RL������\�2�2eU?A�Ѐ-�v9�_��x���U������֮]%+%���ׇMD13���>�Z@/�v7���I�,P�&���z�V�N@hRQ�j ��C!��IT�3�r�SA�%$$�
l�]���Ⱥ�����g��6������4KJJ���$Fį���<�LWy�K�{��Z+�U��g�ASb5S���C��5��]\���_$���Ƣ���oW8cg��I;�ځ���q�F"���^��F%�̘%Ւ�@���Fb����la����#h���8�Ի�ǥ��tw��i��V��ۅj.46:��HkίVUSc�\��>ϝe�g�;��V������C�S!�W�36�-/W}��k���ں�𣝍͚��e,1r� U�}��ܭ_�Z3>��/���!�7���f�OJ�@��XKB���ۦ.^Ak�n��*Ea9(��0��@^YzI\��ד�5՝�Ÿ����.�l40-n��D��΄:V�+Zy���J��<���=���%Ѽ��{3>��۲���T�x?��º�͖E�5[�4>���A��(!@�Xߣ͞��ƺ�tȺ+_v��^}�����)M�~s�����������N��A��q&[���q��Q�����z	a��6�#"&��]�3��RR�o�Պ.x��򔕕AP�^��?�oj��a�Nc,�������[D"ꆁ�˕����m||�
���ޝ�kPmVʓ������0uܴGq�θ���u�Xdf���m��!w�af��ե���յ��;�i���؋�rW���J(��~���/ g� �o�F�4�p�%ԕ�Sv�@�ڿ��n �xP@"!�����0��������R�C@�#��~���un�jP���b��B;ŏ;ac� t>��}f�ûjN�����%-J+�4��MiX�5��/^���z��H��5��H�y��9�~���9 ���m������!���2�ňS��w���z�����U@���70)�����;5!�5b�����/ܣ���d�c� ��=�>{���L����ؔf(������ö���۰���j1���0���+��v]t�E7���^tQ�9G���v����`f��&%3�b�'��(���I;gz��%'���;�lG�;2�R%�neiy���A�*;fw�X�i��C���*b*L��s("����w���*o����p4�ˈkD''�n޼yd~�VR]�� �3s�G�d���f�;��w��s~�j�lr�m��R����幣3�!��6|��4�d}�=�!j¦|f=Z��Q���܊�Jzi{��,�0XҤ�=�,��*���&A��@P	8�Sm�樺*��,�!YYv�RY��[�A$$'���ﶼ 9U%��w���j��>�0���̙3�(�w,�<[`W��$������I)��n��F�M<	2�xÑF��yx�}q���/}I~���H���S-Q�c�dz�}��c�xTQ��fq�E�ҚW�O�yxx@�Ƚ��R�$�?u��4���nԌ�Oj}k�J����ؠ�z�{W�#������%S��n�ef璳�D:�OJ����ȞN�h�\3^�u�\�p·UIj�R5��5��8�0U�'~����ŷ���X۽�_Ks�a�y����e���+��6���b������ 	����L:\~;5����q�:��� lh]3�s�%�����\��sL�b�W��-�G�lه+���V���W�aMT�U�eee�~��n�vO @����t�bAl
�;%--va�����`%�Z)f��!efB3�x|��������\�`�xLC��k�F=pލ��yK��}0�M��w�&6_�k�.J3V7�y@O@�.�]����dM��UO3|�[�mL���E�<�11���IaD	��ĉ	gy�)M/���\R����j�֒Vl���rr`(CorIu�� H���^Ywڣ�~��C���Ffн[����1�,z��f>��\�H�kmy�'�}*-��km� �œ��,�ܮ�a����ځy;�#��ݪ���C�#B���<b_*=���P���]~���đ�y4��ť���oc���_�|����D���2�&O+��XND�|�p!�O�x�B���!%�Y,�R|����m۾�[�z/�����Dܩ���!�\H{��5 bw�Fww���y�:��F� @8�F���\�^@�����VO\?5��WTTt{����nPM[ZZ�Ú�3��a����-L�L���F�٥ϟrL�G��iՠ0Ndt4�.+����ƥ(?D���L�����X�'�9�h��>�F��f|�c�K[��pn�U9[�����_{{�(��x�f�	#�]��p�q�(O���(����-�Ġ&,
F8���v&贠�a��I�>U���:]QQA�&?�ۮ����T�%��_r��ذcr-b���Ձ�����m��O��	]0600���f���NpeЃ՗u�n݊���x����)�v+�Zl�������ݏ���V��/�5���M6|���l�/��"ɸ�ש��Qc�����g��D�+�Ū/�񞅀?�@�k���E��*u����˻��J�/[�Soѭ�-B"Xu+����%������ ��2Q�� ӵ"�}nB?5���⒏uS�`����"���D�O�>c� �D��R�%Q��z�0�_u�J�yi`$�a~�m������f�;M�FyP�h�����R�i����<vw��Z���i���r�G�F����.��&�H̿�6�AiS��CQ��:��A��6�}Z�v�"�|�B#!SAA��1��|��~=��#��0�dC@�s��5f�gⲟ�Z����{�#�_췻Vcna1��QS��P�`�ao(@��gς�֋��EG���i@E�P��zjٟ[k���>�x��e�<|�[��B�P�x���ZQθߴ�!��@x��B�R��|s�L��\�t`����:w� R�u��|�O<~v ���w^��Q+�y�^K,�?X��.H�X?���߹}���ᎊ��Iz��_-lH9� ��vb́{%��^\�&<�A��-�lW`k���9���U�ς�EyjtO��ǈ7��� ��h_�iB�kLj���1�������6@���'A���Q������z���3�{_Je�DF�s#�jvR> (�M�"}��)� ���:������R(��*��X��;�)T<a��Dǆ��"�ب&�:zݬ������!��*�	O�{��䊧uO�8&�7U����ڢ)Ǽ�v4|�p��n9�r����ߙ���tI52=�t�#����缙)ͦٛ�-��X�����t�QC���w~��N?� o��sxX(�b_P�_W���2����;�m��� ��|*Sq�ż����7���U(�kg\T�
�o��m+�ۘ�����,�_�F3���<T��Va�Q��6�����0��]zv�cE����t}~�
0�U~��׽�tW�>�=�d��J����U��q�������3�`�O���b�?r"(��|�ԉ�����L�S�G3b[�`�h�d�KFԽ~}�2���eT��A�U�}�����Hœd�h�D���1�I&��!ۺ{�cn��[�t<�7�&��N�s���Ȯ�3�k�CtO��"�@H�6>�)0���4`��(�ł[�]#4��oڄ�b�D�����<s9E
 ��W<�%�T�����<�K*�,��1P��&1�Ɣx��8X>Sm����h �|%�{f�(��,p��w-�XB��'H�,d���QR�7��&c�W�s:�rnf@Gķ�Q�^���_����5��k��
���[wP*�o�GM�%P5���C���M�<�"M�پy�D�5��`P�{��EO$#fz"���L�p���z�������B�}N��x�;��i�<l��v>����1GE��[}�x�֎хm� %���?��׺��C��RLtS�Ⱥ��;w�خ��y�X�+{�ej*���۴�s���ձK0Rh	}�X����һ���w�D�$�6��I1��xg�ndh�*����0�*�y�τ���~�_�{�	���g�'��O���G��H_ﱩhO�KY3���'ǀ��@ �H���}JPޖ�b9�*hH	x�1|Ow_<�@�B�����x(B�������޽�u��Z����I�c�����A��������+��5���m���#��沨��;�f�<Z��g���x�_X�-u'[t�R/�z��y���l�Ak��χ�Q���(�{��	����@�֞���c!��s7U�k0��qʳ�8�Iu �1Yg[�޽�0=�?��n��/�[2Wc��;�f�֕���F�K�v��d���Ok���Xv�M�P��\<����)��@G����d��iŵ|
�L䙬P���NG44�3�=���Ԥ|�3��3�:m��o�~�UBB�es{'�����Ŗ�Nc]@�$ �M����4F%��=�m�M���DA���&_��پ���7��d3�fh�x��]��>��n��]ml��M�"T�����ެ�F�//�(�b��u���L��� ~���J���+�#�r���[JH�����/�i��&x_>P�R�;DK�Z���hhr{���<�%��B�(>��3]#����HMFk��%�����}Un.�1Z=�O��w�lS��4�B7'�O]��d(����-��.���s$�[�@����7�B����1�@	Oi�h$�c��f(å�R��k��>"xr;�dʜ�ԕP�%���R��%n�8�2��H� ���a��];4D�v����HEEe�{
b����j'�V榒"�(-�M�dϿR���kh 2ǯp�jQ�G�z5�������'������$������=��D2O�G'��߿��s�(C)��g3m%A{ݦ>�N��zؐJ��聉��v�B) C">�� ����u�B<���]��,f���:��ŝt���$�X��ϭ�)3&
a�b0T
��쥑�B�bB(�@L�i<3�	��T���@+/�mfR��I?�h,���{���*��-�z�mO��h̛U�d��%/��6r����8�>֋{��q~����5�O�����^�hȕ0�����d.?KXQ��N�H����� ��5��_�ڐ@� ~
����$,�@Ծ��p���-�`t�e��̫��>F�	Q��B[<<�ݩ�*�ljz=���e|�/��K��#��[A���;��K�w0����d/��_�@%�_L6�����:���� #1����T��l>�C��6��^L,�Xt�c����n.��k?���
�!Ћ�\���U�۫��W��|�
��|Ƿ�vW�ܚ�l|�L�hH�Z`�P�SWs��U�6��)3�d�;"5�v�hyy9���Q@�*T���#� q�����V�O�f�����훆�n�@��������"��<I��e�ԔaхꙁS%�����q��gC���!��BހR��R���].Z��'����NS�˽��S����X���51��@��U�de=�����EFFb�2�)���������.�AڸriK�
J\�.�А��K�{�L=l&�%� �tn=zLU �s�YT�k�怐��*�/ �[V�I�P�#�?-��S�2�Q�f8			�^_ҫ��鱣q�M�8�m��aˍT�G�Fs  Bи8;;�&B�22�i��Tz��������� X�hwvpp�.��>ӷjhn���-�#�DṶb{w�<,�f���ph�ݍ�N��1W0�-�f.�ӹ�����v/���x��I~���g<�~n�9�#�CW����4��UK������UqkxE�U�u��ԭLM��\m� �
��+�iX��d��`�>H��K�`��?D4Uƈ��1���`���|�-f6�����e���!�'!�Nm�Em�|���~���3��@𼽗���칾�M�DN��U��2g(\r�L
x[f;	@���?��= 7*�s)i�::��knHYZQY�/�jL�L�M�7 xTTT�nv�=F���P��3c\��F].�ı�<"1}�͐�C�%q�U�sK�P�A]�?k��ܝ�X����?��#;���bm�w6&뫸��{�h��

/>~O46q��P�ݕ�f���-��T�;����3�D��T�*�rN�};��&�V��$˾˄��Y�p����DW�z�[WRRZ�=��t;��L|KK�������Y1����|>�ń�U���i`�Z?�Bu#t!�v�L���WI(���-/<��O55s�5���� ��XG@���p�ډ]���h2?\���˭
91޻�\ ��k߃Z��B�P>�98�HQ֋ET�>�r�W��y8N?	�(�ĖI�g�����W�gK���cBS�Z�z���,���l�^k��9B��u܌�7�>�={�=�u1/r���3k�Ua"��(�|��� ��''��yϚU�I>Ae�J�@y#<^?Vs����;B�=��&�NpX�I����nXoffv�kL��%0�(���6a[v>�a 9���yCf��E"�)��`7�f]�$�]�٦ŭ�֠Ya_��o�%'51��؊J� � #����nY&&&ݯ./�s�n=�h�t���<:<��a�r�_�v%�s###�<|C�^4d�u��6�Zzz�V��{ѴCx=TX-B�n�-�l5�T��u0a&XQ���yLNf�:�U��VA�WEd�HNps
7��Sm�P�[ʢU��gH
^�&�T[n��BLCm�n{�sZ���X�����RJ�@�Q^#�����B�쭢dD���_����x~��޾��N�U�f�'�X"k��B��Ԓ�?zNZ=��=��'&�� "��+ٍ�yѲǵ
Y��"^�0��������Swq&$Yd� ��)@���'�'!]H�����i�B!w�ݣT �僄Y�Np�������q�΀�X�J>B'��n��<4hO��˻M����Y3�Ft�gY��6f�HJ�����aZL�?b�7������C�&�: |�K����/���.��v�=��bD����
J���ǨIoz9�+�<سn=�Ye��r���lvlvZ�t�e�5�Z�O�����L�V�����]5�<а���p�&����	��R�X�޽{�sc]�Gkk��z����=]]����(���/P��D����?�d����db��J1� Xb8ɠ[Yщ����i�U��GZ|;�����?a�'��E�/�j�*��)s�������έ^>8d��X�m�����V����5�[wb��kk��YYY!�Dy���pe?�QQW9Mc;?�H��A�`����`������a�TS����C�P�ц���b��P9�,L ���S�=;�)�DwRy��ʻ'v��0wl���#PӽU1@)��"ؑ�7�#���K�s��K�.zz��d�>\L����ˍ
�V����tP��_u=�m�77�	����/��;g,[d|����и=(�w�����i�DN��)l8,���NM�;�<K,�nG84�V�Mn����-Je���A5�)�Q�׿��LNN�/|���no�g�2z9��}� DcYj}7:t�F ˿��q:;��� �<�n4�~=��|0� ���6�n�V��봰6��k�9k���4���\2Z�=|��Y:F>/�r�2J����T� o��%k	� G��MXweT���lƘ�@�V�C����C'o�!�u+�Kp@!�O�Q���2����m���]>�OXX�u�$������=8Ce���Р>+Q#F}��[l�C3�c�wo%~b+��O����L�"�v�<����:��/uA{�E����$���y_x��ꨗ����?Z���7;�bqk{�奥W����+�AN��U����j���[>\>��ȓf�K�}���Iw�����!=㶮�'-��s~��H�2�qv�Q&;f�9���A�*:��_��?�1��ۻ�+�>���3��A[�JbMi����8����Zb�Ű [�vOV>�jA26p���o�q� 9�Kk��핳�_�ĳ�g��uSܗ&�R7J�5�2�_���A���*�E�.?d��9�m��5�1rAΨ*�����ቭc�������;'v�ϓT����B3��"�S#��i�P����@n�����q
oNC��a�zdݕuk��ⴸ����z�V-�����}Z����!��.M��W���P8��dV⭩Ke��YCé��������ު	T���{�` ��`�d�k(V�|�"�2�c��o$��=E��o�=�X����U֮#����7�U�Z�}�Ү��$�~�M�T�f�������0����dts){�f�)a-���� W��"�����\W�����4�u�zu�;MMA�}��2������v��t��\�>#L�N�1�!Ԙp3��.���c_�*���P�aMbU���WTU%a�>��H���'�r��E�8���:bb�2�߱�1XM\��)@k�q�X����/��q��JC�8`��'R�󟣫]���I��>~��d�Л!�{�k��[;�����ˠt��(��H��x�K���	�\�<~�Gx4�A �\]>�ߥx`� �wT��@��Re�%���6.9��O��vx�����O��ʋ"�i��}��l�V�]/��$����]?���A >��޾��o`0��<���+���͍��w�$'�$�m�Be�_Y���/��,<�^��i�GY~FX���G��_;��-<З�k�~)�'���T��@Y-�2�Pk��)�Jt�	z��X��\�����wa��*��d�Y]�x�{������OK<m.] ��/#`u� x��ټ��7u�ఓ4��c����"o){�5X��a�v����yx��>�����4�b�_�{^Tt�����Jv�Ganx�CzF$��Q�6*3�X[�:Z1j���@��p���w>Ʈ@ȠE���f�z��s�	R�G�'�Ĳt�U�X�R�{&�ߛ��l����S�ј �_����!t;���y=t�p��j����x q ���ڵ���.��p�I�?;5���*�8&V,]��1X9|���q �c��p���R5C�#\Q;��L���Fn�qOv��i�<x��vAI`����G��� P�6�����N�i�A:�آ>1�v���h�Ž�e���^&''�9\8���~��QNǲ�{K��^w�ݼ���ތ\���>������m4�*F���4þ�I}ߢ��*%t��\����]�{��QJ!��G�5�d���o�'���n��)����>�z��R�����o}��K��5km�[^4��]Q�8w'���<r�����-�<���5�*�����*񓉿`{�x���}�v�������8�w�#C�`�g�����8�HUαM��s3)od�L�\z��ʓ����pF�T?��kn�v���"""�\�l���i��'Ŏ6����m77wZ4���j��=�\+����Tu�D:�Mks�.����giF�y�t�@�u���y%�S���M�	���_H�Mݙ��W�v��Pi*?M�ƞ�D�au�5Y'P��w��Br���X	������q�"�^/�u�~�9]N�BU����o�W�Pu@�C-�������5o˟XE��v=ټ�������^ǻ�qǢ�ϑukN����V���1ڢ��6�>�y��h����YKb�h��������R�+�Ŷ��j�#|�Rvm]��<f�0���}�*�����yA=��a#�2�7����������뿱���!җ��M����Cs^���z����T�]������,՜+l��C�y��D��!���300�@wܿ퇉���9,��L���m������'1BMH�l���]v�a�uB��Ύ�O�>f�����Ox���Ii���))zIu���pZ�, u�TH�Tz�j;�%%� ��^�Z�����?I�˝uLw���2՛��3	w�� ��w��y)�fo��Q�^�x�3��~�a���i��6['�#3�$��d�����̙^�<y-���4C�]��+��H�#J�N���)�9xpo&�]�=�N�Lo������
MMۧv���=��+����+r���K�$6��v��1V�a]ۈJ/L��j�6�G�;p5���C�c�c����&��%-iN�&GF~$�9��@`�s����orH))&��B��3�9�Ƴ���_*�~A�a�����8���m�N���X���7r��hIV�|�9�����u�U��m��M��ʡ�y�1U>�9�k�(P�/v��v��6���I�"Β��,U{�帏����0��K2h%��ma�{͎��M�x1 wz�d�6�*��Luh���)���yg�����L�*\���{� �efK���!��w�2E��X: 0��
-���'�����kHs�jD�WO��<)� �a�M�E��G7`��R�ߏ?�|�K?)dĹQ^OLU�&zU^��a�����=�a������/ճ���`��xq���b<?����TJn���Z	;��hp���C7R���G���8�M�zބ��w�~LM-�$P�������\���b��{@r(a�|����K��yŜ��#�U/C��Ƈ �$�O��	�lZ� )�ݖMt�v,e�03ҫK(�TOWO�GA�^��L���!ef��2���P0ˉ�@h=mnBL$�l��DC'f&�8��W�Oo�{s�W�����Z|g��3Z�A@�ec��]䕥2lоV�������8�Bm_ѐf�G�$�����Dc�����9WB������F�Xt[��ޓ8Ҋ�ɬ�{����L\�(a[mB#��;@�?~��=x�3�9�D��ȰJ�ղn��SA%�SM:]-�j��5��P���6X�n�U���Yv3W�,�3�k�sg���s�_�R��T�)���(�F�1�fB7�O֌YWT�r%���e�y���y���r�R�C���'���mG�>c8�[N��4�<�$����i�[�@e�Y?	�A�֮�q-��zM}.�RC+����k	Dcn��$Q#�����f��Բ��dMؿ9�(�v�K�̾*O3'5ѝ�K�'���NW���f��У.�YrYB����ܻ��{`.�+j�{�u��Mt�XX�r���t鑤͓�|��G��1���4�&�ߋ4JNpncd��j�p��@E��m��S�mo����ڦ���9{y�T���� � �'P�HF�f��=�a�'s�0cA�3��x��f���CRBܴAZ�AJ�Y󃰐Uԋ�)��÷��05�$�Ct�&x?&7�/��J�4F��rUc`2����ڭ�X���|���I��2�������,��vZ����׭3[�4⻂JL�&���h)��\?~��aۤ��iُ!�IX����L#R��H�F'�'���g����E���o~B��Zq�3��m~����C�����> ��������Ig�Hs̅7�Yt}Pa�-����1|���Le��������d�efp��C�����h��_��$Y��������V&Q�:��k�@�FN.i���C�$�޽���u��b�7�w��+��y���{��_�]D�Dcb¹-��^�M����0�h��y�$#2K_��13c��gX{A�Z����[հH,+�����7&����IL/��������H�W��J��1#Q>y������z�bE�����juW���4R2z
0z���R��ϿrH|Q��Ƣc���V�D7�XQ�]>�@����-�Z�a~s��1�[��7V[K
�#ď\5�����
!�{�L>T<h[Ĵn4��	����<|��Z���-��P�m>��C�'v�p�NJby(B�����!�B��L��b����p�`0�L"NQ�������t�^O���)��*�c��h.�V|�e������D[X��s6`O�.T � lۣ
U�ŭny�Oo�i�7D��v�:�옷(�������v��s�s,���c�6��ل ���x͝���$���[]���i&�Yn80�QD�Ɍ��	�~"�j2���HꙕC�����(�$�7?�X
@�1�b�[tr�n]	bq����l�t��BU��/�(Þ�c')¼�]����	�p�/t/_�L_�sn��T;L�^G�>Ļ��8R&&�gQ􅥺���6ޔC��ڞ�hd!��G6�F���(�h`��]4��@4_�YJ��ѿ��E��!��k���%~ q�Aa.F=�2R��6s����G�����ڷ՝S��L�!��Q
��'���9��r`�my�&��v��z��e�{��&R�.����
�7����&�޹Ô��=z���
46����@O�
��.Ԩ��l����"D�0�U<��w߷Y�����$�m	�a\q��QM����L��)x�O�`	��B!���ؓɤ�i�<�1�a�c˒��߅����t��;e/P	��.�c=�*H)�"��
jf���:�f�A�d)$&��L�m
��G�z�/{��۠�fy���=�6O���p��qH1:%�6|wV�77uQnL����"3Ӯ��NuAN�{W�x5�k��0�v�|O��꜊�PV
�su·�`�s�\�3�~�k��95�M�9�H��?,���wwY��%�'�@m_��b1=4���!����h��Xo��8#�~��� ^�
��`�jeG�0��h�/�) �FTD
d48�Y����dZn@|�m�_����A4�΄[�����5oNj�u=b��� 6�e� 蕰<W��73�3cU�	�0m�&Q#�(Pl��[s�����0c�J�n����v}<S�%vY�+�����󇣘3\�G���D8s�����D{��_+6-��=#zg  ��PN(�lԧjL}nX!�$�[^4Pw�d��²���3�ݾȡ�by����@Q�'[^@��A�,gXx������-Df��kk�P�/ac��k����Q�-�YW�l��->S�O
Rp�$�s���R��֏�"�*�A_�h��͌�&]G��57�8B�ω��v�z?�����@E��2z�P����Q����YZ�8$��n��ͫ��^BwYh��U9�y~0��K���	�,5?l��|�?�M���:�rTE$�6��Sv؊G��<g6llC+�K���W����de�Un,����@%~U��0���������/�Q�m�������:�O�?�b�b�O��rL�ｔX;f�|l�������@3��C�a����G堟��zhl/pfd6�LL@��V�\�d-Y����_fl�ņ��Q�yltX�Rֱv��le�$@>7���n��E�L]�Kגd���>8���^���؆^MN�(X����kW����B��5�B)Z�u[����4ڴ̴IHBj��2�$�1ej����&-ӪFj�֩���=gr�Ͻ�{�9�����]�������sLJ��"��4�|F�����gjh'�x5E��K0/��8A�`���,��!]��;�|q�+�7��<L�-�>�A�b�h��IZ:-ۭG+���u��0�D)��C�Q�&��+Zא�W}�okk����w�IAHi��B=�Y�X�����A�xMwq%I�2���o�$�*�$��A=ݪ	j�:#�l]T�'WQ�m����.x|<���L��������W�Cci�w��Kx�QbE��;�o��pJ1b+^I��{T�^���,���	��:�<A�yF��"��P��<$�eB�"X���=ɡ��ml<���'P�����Lh��il$Y�Tf�P
��C������{��Q�-q|��6�^��xR�c�]�&�W�lW��ũ![�����%8M���aE2N�Qf����ݺr$��OY׍��,V�(�h3��Ҕ��_@kTu��T�"��PW��T/j ��o�ow��֏z�T+�bZRK�C��#�gtY)���m������{����q�jެ&D��1
7i�Rى����9=�.�K�ܑg}�|��rf";l"��pz�P_��
=�����TÎ��WG)�K<���gp����ռ��H-k��ϺȚ�n�`FN�SY��ůۈj��8���>$��p�����׺��39H������5ԯ�/ V HRX2�t@���S�j�o:�~����P�-�҄�~��F�_5-~Gz�uF� �h5�2����눴/���Bj�6$�"��ދ�VP� *��-�r<����y�~P��<˝�d_��	)ӡ%^��[�7��Dˢ����͌DÄ�U6H��w<Rp �YD�h��
I Z���u=��I�
KZ�I�ۀ�Hĵ�wȀY�Q����h��R
���Kcd�HIIi�� `R�^Q��啄L���n�0�%5g��d���R>3z�`��8�Z&��+����"HD����gQ�n�n�!��e	�7�x��y�F��ӈ�s�:�܍q�ׅO�d�1>� ���<�!gK�͔C��#�u���0�!}�U�v��L�����>?Y��r��rVU��'d�4�ƌpc�­�C�]hY�o������#k���U�T�g����.q#��X��g~�s���2I�vm�!/��f�v�V�[H7D��n�k|~C��4~�jw~���ˆ�󝕽�2h	�ɀE	���GѢ���}�s��0�/u�F��L,\�J1X^7����Ul���C\��m�QUi�����tVR�͓�q�b����Lh�2��yl+R���ejBG�)0\Z�����Hҡ:Dg�״tݤ(�вaTVK�JН����A�O����<��0����0�����ܢA� o�L�,�����u���s+G͔;ۢ
��?�Pʋ������#Oٚ�$;C.���6L�zt{i�����y��˵(*|Ӕ��B�w ��+M���
�$UeG_���t�ؚ<�U�	쑠��*��� J=|Od��[�I��N_
_v\}Uf�`Lﮗ�2�ed��\X,Vo���փHi�ؕQxB\1 TA�#���;ri~��RZ�wv�c��NP��{��+���:�N�M��fn�Q1��0��MhMK
��O�Jn((�8k_�up��~��^���������f\�J��G@�re�L.	��17�2����hB���lP{�?8V ��bK��3��짼�Qt�(�V����dUݏ"�<2%P�'��%�73-n�C�W'�$�����0W��;�մ�tAXY`�R�>�
Xw��\�D>�+�:)ʊP��<�2+ `���ڐ]�#�����(9�
����q3��/�@EI��z��)eeh�	�a�ܢ	�Vâ�B��ىG6�K��(n*�0/�/*̣,"k��C�ޗ�����u[���ӔTӤ��>7�6�}i0%E�zSH�3� �f��Rs�]�_mG6���>N��**D92�4#rme��}lH�GV}���Ɂ� ��Q�V��s�$��~em0tHE�Yyx�9YLg�0k��z-������`��u�V�\l����p��s?���Ɣm��v<)�~}�Ŵ��st�@mKΝ����"�\�ʎ>S�4p�2م�����|�bA VuA�7��~��.��B_�B�w�T�����_2?�h�NY�ƪ)���[���_c��;?� n]�2pnm����V��LQA���3&3��f�͚��͹o����o���Y���ە�X��n�XQ�XP*�·xAx���e謮N �'�G��s����O�T.�Q�2V����++��ؑEu�	f���C� Ȕ��	��'d@n^2�* �U%fI&��M�Y��y鏏f���x�ѣm)=@ ��Y\�M�����g���?CA9R� �*Q�sA(��I��{�N��77����q����I���ć�D?H����$��)�h�D����Q%~!���C�Q�J������H�+�{h�� ��t�5ٔϫ�`Ƀ-S��ONN����*��B]<xkGD�jef}_��P��t��Qz�m(
D2v�>H��Ǹ�8�	6�7���3�$��(5m[����O��Z�����(����,�ݰ)*�����g^���е����>>�N1;@[/&�[C9\m�j���e�����S)f8Ah���)�w ��(�
Pz�}�ywC�k�Wu�	�������8!�0�������6��,e�b��\��.�|����g%���q*��B�R	��d�>��@VYoR�%V^��3�*��A�694�qA�MҼ�%���Z͍.�vq!�ڟl�P��e��J;	��\pLo
6��6���u�P�����I��@�w�Ϯ��/˛�=�SD����Pq�z��G��{����ܷ-h���s!5"�����9�a��?�rz�c�@8ňn�����7j�ɵ�ؔ �[��E��.t�wf���Ҹt��j�����f�I���1�0�{ ��:Kɨ�bS'�p2��o*uV�D����&j�����t�{��v���m�Ƈ09.Al�ٽ����&��":n���\�n����J}N���GMF^��@��!ڟ�w" bG�;�H���|E�{��k�D0?Rc�����^C�͡K�%��:��yg''&��)7c�4��#�J���R�Y�~���g���oŖ|��� b(د����Ǭ����*r����p͚���;O�2��,y �R���(���?�b�9J�2�e�#�!Hk�2��~��^�V:�����{�;�>?K+Π������Ȁa����	�*JO����_����h=���g9�mU�����a�7O�Y��+E	"I]"����ڡ���
n�k2�����V$K����6`o�״7�^�X��k�"��Ҏ��S�9nn�q*u��ɱUXl�)��Ԅ }����u��>���vc�
[�繞?+	i���iu<�^�t�ڄ��l=�գ͏��G)�r�ҿ�tz_U�l��~�Gř
:��5̧p�$���� �\��НR�}��@��j�l�Nj=�V�iR�i�3?j���B��Ղ�6~��F�ی� �m��q���0�3h=�qĎ>���w���L���Ec��ؙNl�i��ψ5IL�ep��	h�U�|�0+Xw��
;�1�C���$�����Ԫ�`�A^d=*���5�e��~�T���b˒�~�)g�7M��ݔ�p{g��X%�R}�DMg��c�j��^t�x���m��J�.�Z��=��/��J$N�<�k��"e��V��^8ß��&��e�V]-��EcX9u{}��7ى�ѷd���aJbD�ʏ���_A�����	Ʊ!K=��u�or�n20�7�Z�(	�����1@JR�&0�������\A�����P�vT�X�B?�<u�q��}�U7�x|D��g�����)t;dr!5d�&�<U���^z��)�"n�Y��)�5�9��l�+����k��P=$�����)!/�U�`���-��'Wnk)��|��p��+L�8��:\�0hw)�$�φ��9�=�� ��T_�����Q�<�%��r���T�����9D����p�\�{֕iL�t�V�&��rT4��[li܂�<гڷߖ<j�N�+�����q����N�4�ݞZF#���$ vTe�B��~Vx�d�$t��H�-�Ub�
�Q����M��t!�����'̘���f%�4�s:���M���7Ц���^��4G��؎X���Jk��$�ۃ���m�:�s[��쓂�ؤUp4��No{y|�R��,O�P�\��`�S*�&[�%㏻f'�咜��^4�=A���A,9*��*f	���M[˹ҡ���3�.0J�H*�ҙJ{O��.�6��6�^�d�������k3�img��˺����y��?�,vBx
����BV�˽E�A}ׇ��+�O�#=t
~$��tIt���l�+����ꦻhX�_;�����Sߐ߂Z�1Ur��x0@߾$���8��υdU�%��a�D��F�K0���vvT���ԝ�g4HDr��s�y6��G��uUUT9�y��KD�\�S&wmg�� �E�4'�bJ��}��'#�P������<�5����3"?�9�x�Y����xv'�N*���Я�?F��m���T妌��\�:� ؅�)N�%��� ����xň��\�āj�q��u�B�Y �jT���:�9ъ�e�~��V�T��Ր�"�p���ŖVn���I�F���I������9℺m�U���k+i=�� Ќ_��諬Q���Y]�����9��L�,`>�d�y_�e���|T�Hd �x�z4g��@F~b ��"��OvĖ����Q��s���L �e���8��F?q���{'4Y3�r �?�#~�/�`�N~��(��Ӌ`@Π_�)��#ܬ�
Y�o������R�E
��Ub]p��$�Ѧ@iB��\��P�sb e���m�0!��5{!�-S?��81���pU|~��H��UW�-S/�?�4��u���\]����k������5�x⯸pz7�������>����O]g��Z���V�{����GP	��z(��u�Q#��ٔ��4�/�S;-p�3٥'w���u��	P�:�{.U���f�&��=��	ƈF���]�%]�l1~3�'�]����6�c�����>�޳��@ˍ�q�x��b�;��E�Ae�25ի�=
�ՙυ�A�0�p�%z�`�����5ď1�P���z�'�ۈ����i=�.��㫫��nU}*���e����BMP�������4��:��c@��=Y��A6&��e�H1\��p�w;����٥!+�#GЅ�]O(�8w��@($�8��,��@��xָ�X���2)3�:q*I&������h3�W���Gpr#��4n�=����A럂�+��ۜ�9���lquI���,n���M!w��8�>�;��/��sSx	�uKD�h�WV���hT��E!�\$ӥ|�^ऺ��RՃ|����,�d���ɾ^<��{����4'5��)����J)=Z�P�]8�O�����{�İ�x�w���m%�<���Ҭu��Q���TYF'��;�*>0rs�fM,M�������i�����>�ǹ+	�������@=�lh30h�A믛��\ŖӋw��r�����D6ȡHL6`�e��p�1��Lߥ$ӽp����3���@����U��>��1�8����g =�>Z�u�D^]HVJ�"GsL����C�	IF�e��e����XP t�k�4?J���K�8)]˰���#�T6����ޯ�wm۸W��NQ�v�,���?���ܳ�9����)%�n�OA��{�8���eI�'�ڧ�I`e�@S��O>�e�)͎�%i��@���^�>�p�
����9��~ھ��:�z^X4��3�#u��o�C>����� !U.����7�^oRݢ�M払kH~t���+�d5��! 5:<1����z�!�U�U�:l�yM�������`[�!l}�^�DE��,YZ���J�󃛹����0'���ك�O~sx-J��C&@d�a�O�G��`�p&�R}��Q���Z[��7����ꝫ��[��ִ�w��y����w�]��Eb��B��#� v!�,S�����¤r� 9��%{e`�hˋ����K��:�)BfK��-�M���t��9+94?�17eبu��-�uq�gn9��7��ng噴�}��v
;��[��=r��Rrު>ǌ%��E4V���n��u�t�=F�A��R/�ܝ
s��
,	�i���#f�9[��ھ_��z�e��5Gu����6�#m��L=�����H�
Ğ��F�����[g�Jg�i7�T��p�p�VkK�&��j��ߴ���#ძXgO<q��*a�&	�52���jæ�����˔����4x�H������p��K�z��=Б�<�<�7�������>#�X��%W��5L\��:��UK������ȗ+2��r�`�"��"���U�~��p�ls?�5�Ͻ�{�����ɓ� ����q�3p�}z��H��Ƣ%�k�ƇW���_0F�؋��LCټn��<�K��\�����
ŁwEFH�F�2�J�P�c���xv�7f�X,�f���eMKbT����;�����+F��D��#Y�%��t�m=����7k�ȥS���y�)5̧�>�Th��}�ޟ���P����O�7����� �m�ОJj���q�y�ql�ǭXҺ��K�N�����V�Uu���*F o�#j!��4>�{'Wb�V/|U���I�y5�+_ݨ�E_� �B�b�}w�ˤg_��>�藏)�����ΫV��J�>��\����V�	|��Y(��ִ��񴞕=H�����r��ִ����6�&Y:#o�X��5�z���s�n&PM|�E��p�R�yb?g�2A��4$��1\$�AW��\�:���{7G�wU�(V��=*�D���\����@T��IX-����	B��2^q	Cf�A8R�8��"qj�����|�2�!AAi�	�S�N�E����O��0�s�k��!L���4��B����LOW9�]��<�j��)�^핍<5Z`B_��H(=�2�î:˧ǎ���JF�m���u�қ=	��};���Px��d�]��X�q "H1��%'+C�5�{2o���fHY:
��S���u��X�����a�Z�)�/	,t����݂?����/q�J�T��X^��듑7CQ:t���#��y�S�
�M6�b�l|1�w�9Ã�ާ��tI�A�U�ꈂ�F�3e�3z_N �W�`V�·��'��3n�{�}v�&���C44 ��#��P�vW�
d���˽x�����5�z��Ͻ��,@���7�X:����J�*u"p�S�t��!�Mk����Xx����%S����X���d���`I̓��ȉŖ��t?����o�J�:<��2.`=�V�����|�ҊsHd�p�� �kv��=��q�冊r�Q
�V���Q�/y
�o�O�	��k���Z��H����C]>u�s'�0�J,���l���,v�
�u�J���Q�=^ڴ(�O]�M��:����+�0y~��2����Y�$��6G���aH4Me����z�V{����3�u?���܌8q�����J�"������⦐�G�׾�G��5�..���eǷ��6�w_ǒn�v;�����u[��`��'d�m\-��sE,h�E�Y�rB��'��=_���@$R�l�mpnt��Ulil�؈���ν�H�/���	��̴o�=16�&������df�ңµ��ҋV�#坨�n�UK���x�����+RXn�j��a���q�Q�0-*�����.�f����h0�K*[�
��ŷ:&z>%w�7�-:G�J=Ƈi\��.~���"
A��8�vJc�]u�uc�RAn�c�V��K3��9��B���ߐ��{���ϴg��<��u��Tk�\چ��q���VǕ^e�5�/�Q�����K�e���2���^��s{��"M�p�,sO͚I}C/�2	%=�o�t3xn|D�u�/�ۯ�>X�|���g4m#b\sL'�\C�IeG_Z���NYm�Y;��������J����e�X����� D��w�e�g N���V�X���^��ye�;g���Pw~}��j�R���R�(��-n�H�"����J���π������G��CD���2@�|p�1��Y��׋i5'�tfH��r��֡:ē���x=w5�	2���^a��q����
\o�
ը(�4����ȅ����
��u*�"�o��!�\��򛁫r�࿅?�T�uF�W&�ͪ�7IL����n����`/d��9p��L�KS����$F(�U���@�6�`�1�iJ�Th0+�z�n��3@~����K�=�ߊOԬ'/g�& ��B"f��|Hݿ�7aZO[.f"���h[y��lB�x	)�ꔠË���E:�X };�X�����s�Tlu\�>����b���<2��L�[��9��$�,s��=!�� �HR);q����ؑMe时ܭl��0qy���j��������wHVAC�;�*��3��UF_�3�����>�����s��$�j6�T�죑�"�$�A��Q������2>.R�٤�{пI�[#��B�Y����V0/�v���nCۉ�AB����� /%;�}[*�BkA`�e�+�NPS_�j�RcA���r���WNK@<�'I�!Зo�N_SSͺ�tu���&���@�Ȍ�vdnJc��^����_��?�[d�,�y]>�ħO6M�2Ȉ��Wʛ�F�X�_f.�@$�o��x�}<��0���󲀤.uI�"��/�p{|n��2�%$�����S*'��$G�'��s����%��aNfk�-�4�=.P�'�j�F��!7��{ŪĞ`�2�7e����~r�a��!5g��=U�Lm$"<}<�=2̼�=��d�$Њ-���9b;�{D'���γL��I4MҊO�ۜi�V�A��&ܱ�C���-��U�5�%�
�vH��W��
$�����F@���7}0#����`� `޵*�C"*F�:���.[$We���w�#œо/uu��<��B����t���	������=�~��@��%9F\��<Ͽ�����Iap��E��8M��,s�w9u���_ܠ��$�A˰Z׀ŐI�L݅e�9���ݳ���N4E�+<�{,��k�jͤ���'iޖ��!��'*D��y	a"���H̯q�0X��"�|�+��q��Yǌ���	���G�<�$d����mk�����?�Ѹ���a5{8�\�)if���k�_Nѵh�:PF6��w^�<�(��Gk!���Ʋ�8��܆������b~�x䢚L�D���Q�r�P|j��:q��kBu ��з��s���b�Ě۟��&���)�MB�Uvㄝ���/�S�a�����@`�j`e�T�M9� C�Jp̼�Y��PS$\�A&�j|b����Z[��+Ig�O��`���B��s���|.N�
�h��z����S�h��Ye�i1��?�/�N��Q�^j�b��딖�ִ���GY�^���3�*��1a�Fp��: �C�bA����-0��Q9iuZΝܐ��2ޑ���<�=���q�jS����V"��	����=���F1�^�+��W'��ݥx��|����Q��@7X�W�v���Z&DV\�J��kr��5ή�e�4�n������n���]j2�����}�I츔����G�3��	<�=ئ>�(�zT7/�jfs��u��ߦu(������<u���bľ
C����h� ]iR|>��Z�b E��%9�M�,l	}VH�>?pRk��`}7�g���`��T�ˏ#���2c�j�r�
[���{�Z��b��>rFM��4��)�V�t���,��Q'��}�� �'X8����2d����}87C$��1��h�L���f"=�Ey)\L��QlyL����s̓��f�]��Y��c��o}���
��l����r��l�-�|���agN�%�J���Y��֒�w�WL"�ʄ���C�-#R1\s�����������ak�Z����xĊ]�X��pe��2O���B;�\L��	��7��v]ǶR�A�Nh�qB�S�g9���D�*�w$<PO�+q}������x��S�c�N^7Y!L?�Ɗ�kn�q}��se��N_l�>��$�P[=�]?$��b���##z07�,�#��d�]�ڜ�W��j2�}�k���;ac󐧴\ ���5��R�����PË�*�OM��#��i'��:��}����X�ܛj@����W�)��%ղ
?U?	_�*/D��}��ed�&n��Y��4mEۚ�˗WbI�I&N�ԇ�$Ӕ�L���B:7���ZBab>��������%�4�*e/������q'��[V��?G��,�y���}�*)���v�l���MC�t�ܶ{M"m��H˰�mc'����O�ұG4���ٖ���f��A��@�+A�p��#���C�$K&�}j[��|�4	g�O���z�,O�s��N�Qz�=u/\�b����=�w��P��4��g�g7���Qz�j�8n�	ͻ�3��$zȅ̺U|f�j�X�~X���'3���e�}>"��u�#4�Y�f��㋴�/_��r3�e�w?��aa���1SY,w|-V�[R^S-�lPP������j݊GVI���S�R��j�͉e13v�r�:;��4�71�,�`fCO1��C[��2I���������mBoa�m���R��Bu��f1/��C�+!P�����aA)����!������k���G.�
_���~����0���!�k�|܀+n�|�,��r*���]u���W����z?����C�0��ۙ)l�X�c��P[KK+�ZlB�9i��yIG�������'v�2�n�2����D��y�9c��Ea��S�3�[d���5��Tמ�ձmd]�OϬr���̨^���V]'�Z�t���%&�EEE�w��=-%e��u��L.^\2�����n��W�o?7�}�Q�����L!v��7 n���S]��Ȕm�I��}��~�}�F��b����5��JO�J���i�Yd�`<мY�36���]aWߡ,?̀R��}{��y��7;r�K#m���}ylfX3;�(nɯ�� ��ҹ
[��I��~�c�������MSRR�;ܽ[����N����7�_3��]�IE�j���
r��@׫)���qx��B,Ľw��w�RO)F�ыJ�1��͛�ҡ,1WA��t����C������T����~�	��p��2g���-4��ؕ7Q��~W�=��|�Z뗳 \l���,E�sد��<��f�R�:;!Z̧�'VJ��Ě$Vfmո
�j&��`��5��1|�T����d�S��,��~��|o����m�qh�����Q�θsh����ǅ��/wk7�w�*��`"K��SE����3*Ȫv �ʧ��Ыx��p��㨻b��5�Fj*�=��-(��e>��ic�(��SfQ���0�m�q��7�&�L���M��\~w�V͓����~>�g���`2^����냅s��7�rX�1�P�h�9����+?��^  ��7��L�N�5^�e}�@��P[�}7ke�G�{/���~p���^#�W{��U�����-��a����(�iZLy�7�a�o�Pg�i�xr���5,���=�ͭ��J��v�(�ybL����E�?-�I���Օe�a�b?	�l��у��3��`FUK��9Tّ-��Fe�[~f-�5gtCVT��,���h����)�3iQ������L��=9EZ���	h��XO�1(/<j�n��/n�r�-�r��8f2��bL�'���}�'K�vm��E�ڵ��Ìyc��t1��;i,�~�� E��d:�2�����`+�H�m�X�7�n��a�T���p�yr�z?��Xr-p�]��$w�aB���U�9�a�ǖ�� �duw��x���<<CU0��e�3��O?�Q���$`�⅚r	RoI�F�#�D�v9YVd*D}��❕��T�Q�������_�7�6��^�8u�`ۻ.N�I���l�aΫ�}��3]�|b�3�F<BuVm_�����(R�ܳ�	`KA��U��@�XL4M0v�h�/����jUԏ�&e���6�������/�~���"VR7��H��dt����uƪU*���rm8�9P��}�m̛x�Y	r�9�O�R�,��7b�7����:���ۗ��|���dm�F��>���{�P.㸥�+�`v�3z6)*�>v�ݭ�=K,3����:���傉NY��s|TK�G���y+JR~�%M�6ZC�뗴�1z�5�0s�7�r%��7��>b��Ev�b	𷫩3�D��7�mhZ��$��&E�%�B� ��,Fx���ђ3�M$�p,�PN3]�h�b(c��V��L����։�s1�Χȵ���}�^�*JNE9KϝF��.lM�|�2g��`���;p�@y�B����@��G,w΂!���V�ny��(������CC��T��	#O�8&UN��:s��Z��'�;l�R�1�Yv3�2,i����Ab����PB}La��$����̆��Ia
��v�Al�߼6��)�u�3�%�_";�\�$��\F��G�V���,��>rєo�$�iҽ����j#܃�� S�1�/;Ny�d;f�e�f&�N0n�	�������/�V��ߧ��͈�����T������������].G﮷Q���0��f�w��i�v�r�B:��oC̶��i9}nS��;o#�0k�$Y�L��%H"�׈D�Ȣ������#��b�=���<���h���'I����3�d��ޠ$�&r0�L��M��u�g�����9?~��Jp��(7b!e��N���EK����T����)�V���Z�&�](^��S߳����>���@9�f�:�D,[�a<�Ŭ�B/�ٶ�L�J��s�=���ց�R��5�3�7�Dh�-ǲ}��է_���O�Z>Q�AQ����lzī���s���̨*���u�'���5gF��7��$��Vl0bs`����Z�bK�JtԜb�(�x1�[7t���<`ȟ�!��c�KMƼ�����sg�%�9o����C���iy}|ӫ�Ҩ��Bk��lIq1�jr��N�I���%�������ғ�eu	�ԐKΝ�靤���g�H��7�9#�̮2	F�S�hX,`�CȞ,�g��U
g��=EqhX���c���r����|�Kq��Xjuuu�� �(x�� �54ߪ���{Y8�{���d���j���;9�D_p{U�
�o�4d�x���ؼW��g��@�`�dC�P�PcqK�ρ�w�ಊ�����t�v�/���R��xl�$�xmQy�'���C�r
=�=�*�	Y�Q����f�� Π�w�N[�Pc�^��$�S��MWՆշ����7��o�::
7�r0�6	���ˊV!��(/ 5n�<����R��.���D�ކ��jY݃�������\P�I&!Zq/F�}�����҈s�,����g��e�~g{��v�ўu����sy�qm06\�Nl��.�@�~�^F5ߏ����I��H`%d�{��qnh8�`��=J�v�Q���o��gx'MQ^�k#�������g���S"/Ci�K�i�|Ts���D���f��%r�Ѕq��򝮦�,LhW��֨G/-�ֲ5����J؁#�!^��o ALy�W���l�����ó��Hf5�?�BU� ���60�[�����i%�N�l4�%����U���xh"��ǎ�|\����I�T��.��1�?H+Σ�cVvUG߹�9�@����=��z��0�����<9ZKDn�9�S7��>�ju>�Z;?pӦMe��Y�<��0��P�0�(������Ͱ��W<�Jvϩ
���oFo,��jD���`����r���2F�[gVHPP�KCU����z?�m�f�=5M�z{�z`AĻN�u����v��{d�n���&Ű���+lAv�S:��y%��(檻�D��@���B��BC�`'x���:� @����v� �^UX8�+�-�#��ذA]f�O�}��O��+��NO[HB,Snx�y]����v��E����c��z��!o\̼�Wv/�=�Bne<���HDzNq�����N�\�E������.�����S����7�[�])[)b���s܏�j~�Q/��Y9��3��9�~������XnKNr��>I�����<K����l���t�b���$-�I����
_���YJ�RǅF	���AdD����Q����m��W Y+� !:������~Ո���Ndɱ�]j�̬ғ��M��{l���-�?���L���jT���iV�QyW�����o��9�~�魉��!j�҈pOU�{c0)�-���<�ɓ'����Z9z���́���r,��\��ķ�zF�-az�Gd#����}�.�rd�9�S�N���W�;����/��x0z�YH�SBv~����	���@��*^� P��\���u�>�����#�:���j��vg��1����J�.�T*0>n�EI�����	�ռ���?�2�J\;w��6nc�{V�������p��1�v��1+f��$�"��&(�t��g��u�)d�1�i��`��SI��0?�Jl0��>/��Ea� ���x�?�m�(��L�|�K�)���{V=�t\�U��W'a;�P:Hݹ�O��������&F㮢Y�;�;�� 8D�e{����Z��j*��Uzpo��*%�}޴I` Ǘ�����=)t�y�BU��O��9�p���B�~��/�=�=�Oڟ�������[O�L��l0����q�wj���1�~	���:����lx��������;�����ŗ�s��d�O��_�1(JIB��b�O���c����M���V��n�l��Ґ�I!��4͊��Ag#�u�׻�)G]I3Mb�r��Ǽ���]��)��-�����龙�E�OY	t���?�k~����
��[����^��%�Ǭ�\jr%ֶ�؄m��'sB�П�{��18����'��*6��w���]��:D�	I�3rW�X��m��s����d����V�P����斺s^i��aC���ȹ��/w{T�t+�Q9)��¸��~�쿩��8�8q��uS$�yO^�9�D��)�׻n�C!�&��l�m��o}l*=��Q��p���)9��Dz'w5�x�ɘ�Fv��,�0M�zZmx��o���ۢ�x5A���o�Q����?�Y$Q҄��͓���\n�e�߲�w�e������DF� �C���WSL�y����~�o��o碰޷l�l����������]����A&��%�*���S�K���fQ��.���ŦMȕ�R�;��>�p����w+F3����k�B�"iD ׏�d��U�w���W�y���E�~ӝu+�X'�#;�R��/�OR,S��\�T[��Y �S�~�?!��I�RX>��a��D���D����@UR��+��a����k��粅}ļm_�yh<R2�Y�%�N���_�;�n�l�߸��Ŋ�w<+�u�b���W�>��ۏ�c�^��kyNY�9��ԿÚP�\mX��`��?���^&zԮ�'���]�Ʒi��_�&���r	���Z�� �ɈW��٪���߭���&_o�rd�z$<	���1+3�Nc�v�{��9)	�)���ǃ�g([hs��Z�k��x�ӏkm_���7���m��|��v{5�UP����:4��yy]"�pEx;�X�Py��rC���bNi�h��<&�<�D�?�.��;|%��_��{8r��/ZY[ �t�{��Y�7�jk�[NL��W��eDC�>E��YƟ(
�Y����z��?��ť�v}�ȿ���*X������3��hm%]��/�%`�P��$��|1&D��(������"j�V�)y�m/t���^��:�����7��g	j�֙e�4�Ջ2E�������{��H�1��\K׶�^1����+a�� �f �����|��5�~Śߑ������#1.����[�� x R���]���ъ
��w����_q�\��aٛD0��ړ�3f��@_�b�җ�  �:�W<����աg<fq�|F�7a�勲� I�pX���*6��T�?Dn�AȌ���
��g�/�}KPF�$p�o|�9�EX�U �l�L�&���o&��be̍v��
�r��!}�C�tެ��Y�n�i���w_�����2�c�htRu�D�\��o��/�"]�	_�Ԗ{��GA\��Ca��� ��m�'ߙ*������`3�)DWl�lR�0�}z��b�����e�1 �Mn�?m�gF\!��_`�or����5L�����_�7��zFq�ػ-�E�:rQ�|1R7Y�T2�}����a>�������������~�z<v/Ť��+Uk�C��2��?Д\d>���v��i�$�"}]�n���S7k)����%��c�ʡ�Aw�o`�*.aF�Тܒ�X|��O��޷�,(��-p#?AϚ�*������!�_�^?�x�#n a�5m��<x�Zk�	kň����I&�&&&w�v�I&�f��)�&��}ͅo>~�?wڤci��h&[�6���HL,�����9^�A�ŝ6��ًo�Ǜh��ęg�.�_�����	U��J�v|92���3�ׯ_��q���N�Yصk��携�젧9�ǝ��_��	J�`6ٟDb
b� 	MdK�YZ�ZH�~LAY�!7��A`�b
��wuw;6/;wF������\+�P*|��Mu��իW?zt�j))���� W=b�Zz��H�������BY�Q����~�z�W;��u�T^���3?>UY�n���#�j��9&���ĵ�x���,j=�}̼	�7p� <BF.ZF���+@D� nW��#G4�ϟ�!?D����(<&�`�j�vjń�!���^������ݴu��Cd���|����KUpo�%g.W��n8f,9�a�{��W���ٟ�?�7�Z����CF� Ba�q����a�j���c$�k���I&'�Y�}L��,��O��8X�����SU��T/���s0w��p8E���ÙX�f�+��ơ(i=��fFuͅ�r�vvz��l9''�qv��UQ�"��Cd��0�_Qq��>��S��w����,�NF�z�m-f�|��e؆5�KHNF���}M�w��������������+�8�gddd^N{�z�LA?���ǢSN`�:���+������zz��S�ڝ���ݻ�~ih��w����I^~�]���a�Vo��DÄ7����Y)x�y5�>��NQ�b���?���ԥ��RE�q��m韃��=E2E�gյ?U��!�R���Y9:"C�����n�޺.C~����J��'zzz�L�_o�:�W���u����P��[o.��AS�K�'�;fD�݋�o��o������M���%��7��r�M��v���rؾ�1W-��v���}x�tYyy�M**내V��*|���W��?��-<����s�����g()��� ��S�f�!��$%������,�]!`+�ֱ����#UW�仞?ZZ{��ZC�h|��]s*9��oCC3��h�3����#_��� ���%�� 1%d�)����ǖm'^C���O脻��̥�+�H��;qv��H@Ӥw�dH�Z�
q	��p����E�G:UUA}3)��͛W'�|ӑ�-k��uކ�̥8x����;��j*���Z5�����0��R\R����>�c��ݬ7���6o^�Ve�sx����������L��E�I�C���ȃb�a13���Qp{a�O�_�[�)/�Ri}{�7�Α����7
[7k��&�F���iО2O\s��h���1�{�\���4�$�s��*����rZ-�����T/z�4$�b/��8U§�ԛ�a������C_Kܟ\���k$��q�R1�B��̮�b�L{�C�a���ޕ)<�od�`|��r�o�:�Z�[[��Ɲ�\H���w�)Vj}sm�&e�[�+������&ih��xx�`vY��nF�陳6u��: $Puʱ��[�{�/Qs7�g�k����Kg�����U@	��i�f�����F������>�&�y��	��� ׻�^W��h���Y#���ط�0�?4t�`��g���̮�)��N���7�����>�L?���n�A�N}��b{��g#�:�����9ͯ��V�GD��n�c&+U^^������#��<��1�W]��^��/�� /L���K2��ӂ,~'�� �J�l�@~��W����1ⶋ�9�Mv <������$�e8I�罸ZM�'/��6��TeuKK���L߅�ՓQ���Z����n��pk�����>��{��f��<$�U�d��kS��W����.c����O��2�m�+a��ۯG������1�G�3=y�a��C��={�Ν��Ŕ���w�`<����W���\x��	3V�V7X��V���[��}�#���>SB]f�S�?����EA���p����	��M���a�AFL��D��U�-o����
�7x��1kB{[0�����U�of C9�w���?��;@7���ܞ+��������Ϸ� V՚Ɩ��ucI�<[	�0 HB�����EQ)$��>�Dqyp�-1Y�g��ћ���#��[mS� T��z�S�]sYB���H�M]�����c��án��qWuE�R�JYs)k�
)BTD�Dd_�eƌ\-�W*���(�2H%Q��B��fb,��9d�u����s�~��u�}>s��>���z���C�J��i�?[��QϬ��^J���,.a=�MӚ�lz� �ނ=nhI���~Q2eE�+8�~ګ~�B����R�˰��=�!VIB��Tq�M�d�D2�Ǭg8[����9yKp2?J �h�Q�����r2ژ��:��n�v���+5\����j+(����m�!єa�ߝn ڐ���Uw�ݾ�Z%�1t�'����랢[�����c��ڋ<{�>�QɐE�<6�jX��d+;;��?�
(3m�K�x����\~��M���PVM����W�5�doyvxk�����R�Ԉ3��[:�1.��%y�5.��oW�	E�Ay���7���W��}~�`~�;7k����!\��!	jQW�|�#G���D2��ܣ� R���Z@�h�|	������:�t���y�s��y�X��%WRJ�p��9�9��+H�K�ȺߐuϝS��"	�'� �����<|��p�Ǉ�R���Q�H.�߇��<u0X��C��&@I�
5=Hm��jH��Q[���/�AF���|e��>�V�9Y���:1�3'�Ո��0���¬�AR�++���-PJm��<���F>d،��B��_���Ă_��-#��t��*.�!�L ڞ�0����;���2i��%��m���-*��r	���?�i�RQ
�H\�pLlS�ϑn�q��ź��1rEL�H@��j��������ɽ�2;i?��8{��:nq�~v��=�����{��a��q`��&q�����4��O�������bf�vxJ�R��]OŶ��,��4B>r�:ɤ�KO�$���q��̞���z�� �IT��7o�J"���4ӫ��2Jg���0@?w�T����J�*��.%�L &fc+=� x����Hi+�4�o�L������N��sX@�1���<Z�����2��S����B�ɻY�F�8��s[>��W�[�~5�{j�w��$>���I�ܰo|�ج�rF��[��[�P�Dq��������*��e��/�XS��D/N��B]��t���+�D\{�9Y�W�t2�t��Ą��1}+W	�k����mఏ�V���.�n���N�h�XgonffY:���69��FMwoj�-ܳ��O��Jۯ
Mo u=�<P�p��Gy���i&�B+w�*���U6_8�1n��U���8@���O�[o d����䪵e�ּ^`Bn�=G�s��Ӽ�eQgY��6a���aV@���sxj@��w.�+�G���������9b_��dO���������ڵ�>}�5=<7K ׳�U�ZH����� �D+��FDx\��G�X���S���9-H�gʊW/��#�#˦&�-r.oo��W��.ʹ��5H�
�7�����S#����>?�S[�v��G�v�r����&��&���	+Fa��=R� r4v�J�jjY �'Y��q�&�UB]��л�H/'D6����9�-6i�~I���n��L��\z��Ț���鑊ѡfi����.�1��,��j	X�be�;nWEHj%���_7���K=-�=�ȡ%۶:l�]������[G��sf�J���BCP�F��^�Mi��+[���Ç������!�~��3&�<J����	lY!az����:�u��GJ(�᷐Sկ<V
z�A����>���EhKA
p&�E�L��`���j��

�v���(�:t
�ŝ����+�
1���:�D�م�V&!h�џ LO��v�X^Ҳ�p$ 3���Syw�7���n�)�LZK谂���b �+..�V�'Towǃ�p$��yQV�X�*p�VK�R�.��pZ4
��IW��2}�U�k���ԀOw7�G�rF�'Z^pBR��O�y�
�T�#�ϝ��Q-ZO;��|8'��S!���<҇h���{[�"aI�^LB�]r^$��e���.G$�g4��ҁU#���!��ȂY�õ<�h�J�QCԔ��	�X����u���y��=*��G\;���h��j~����gϟ 8�D���ocb���[�1�W�čMM��)�xR��]��6�U?�@P͇Bl.0с]_�%�~��&��Z=E�3O:��Ԯ��cG�X�2Oػu���lq��xOXN�cJ��� ���f��J>l���ڐU��9�:{n�]�\�d�I���������WdP��Փv�=(��X�Xh��ћ:ɂ��gf�^Ļ���]DVAU�9@� (��<�>{&���o�$$$�m�vT�p\t��o�:񇹳P�����N3�>lHXTT4[q�'��"���%��@��M�w�0�T��S;�B�U!6 `j�p<�"�V����JN����r
�u!������9b��O�e[C��������p��֬Y3
>@2tu�����e�����0>��˔.G�^����c����Om�<�o���A!S�b����/6�:HVx�:=]���slo��7y(r?�,6j96Y� 	�d��~�	���#��=���Q�۟�GsJ�i�h;��>�[K~��V	��iW�.\��B��mn[\7=�:���{-ÔV����85�yGuu���8�J�N�"2J�4;��CN���@�«�t��3��V\㜅�ߤ���'�u�>N!ԁ�=o9
\��h��z�Y#1C�YI�ɨ�t�5��r(��e1&4���쨌����	o�!�d����䗆�DP"�h4�B��o�Qh{�GT�=1Hu��] r(�I33�ލ�������|���ݗ����ñG��ө����f���S���;�0m���}����7;C�t~�-|ں�rnĖ210M�mr��Sy�k����ݮ�ɨ��Դy�}Y�[Z��ft����\�*}�_w���K���q�}��'�WT-�4��a<�Z�]�q��<���%�J\�}3�؟=��]̧�s
T9���'�
�s�;ʄRÆ���Nz6� w��$E�N<�;���(*�f�*V��yAGK�c�l��*j�uΒ�ι��5��u���%
(�]V:[�x>��hkk�8'\SXQ_�v�=N5�������.�z#�*�fN�%ⴷ����C�r��v���������eio��?^Gmz�}�92ύqK���^~u�ho��hgbj�?���izf��_�}���P���d��9=�CY9����M �j���mV�;.�(�`��|��g�5T�ˏ�l�{ǼQS�"J�����ㅆ�ZrR�#iw����Us�cG{��]*~|@�`��PJ���:���F�E9�C�&�uޅ(��VQ#tۗt�V9�Z�)�\��C���̷��4�͔	���gCC%�L��c����E����`Mg��@�ț//��O����"�7P��b#��N�ww�JKi<����@n��̞B�A�ٻ4��W.��n��"���a�͐_��9���C��C�W[�K"�|���R�� -U 3{�)����1#����ֶ�^��{n�B��:�9Iu��|�ѵ*������_�]48�-|��AXuﻍ�l��ɾ'\�+��#`���ùdr�����ul��_{Fu}�蠬�0:����X�����dv{3���d!��63��|��ݳ��t���_�	�@X
G�8�5����� b2��/��?� ���YYaD�zѮq�̾Ч#��m�S���+_��[h�+\)2�[y��Cһo[�=$��{	����?����T��܄9���]�b|<{�_C�����)W}tm�Q�w�����rZ\%ַo߬,,�T��x�;]���)�*{�Fɭ�UHJU���-|t���Ŵ2���h�I$���Ŷ^��<�@V�'������~	P����ĽÏ Ђ�YB�|SQa9���y��H_ݘq�]�˭�s�@;U�O����l0�;3��[�2�,�z��^�MA�����
���������<9̨�y��k�I����N�g�@� ʽ������t͜����YM�P��<$���'�-��r�2����������Aw&?ޠYHO:��Y.��$�2;���l��s!Hq�5�g~��y޹�҈ TM��glw�Bz[:;X���	��w2�w����G��� ��	#��d�z���VxQ�8��S��{ �l>D�4����ɘ�@����J(����j!��������X˹pR�8�ڡ����{����\H8d�Lk��������Q���{�Gm|�6�j����j�'s�?�H-�˱>'�tn/=4X &G�f�D�@�bPs���nd��)�z�R<�9�)�OF�4�l�x]��J�ֻ�M����C[.G�۝ܴiS�5�8�����$�w�`�V���F����d(TϠĽ���K)�S�#����z�v�V��UA����ΓB2�L���ǒ>�����olT�wTx4ϗ���ւ9��jz4b��ɯ��)u�\�.�C�v1�A/Xh�A���L����11h�g�ubn��QK#��dv����"�۱K�H1�����"�G�1�KA`Ŭ���)�2@A4�5��5��Ќ��@ϓ��"�#\�����?9H$��9��TL���T�G��Q�:^@�D�V�d6�����7�gG#"'k��":73d3:K�EY�3wee��K��0��z�b�Q�]����}��W�7q�S�2]tT0��o�o������A9>���%?~C���#c�f��.��O����o|/neF'Cqs�}nR�#�?y�^���U��5Vg�
hl�w+;��t2R��D�?Z�g���&�2H��j����~�ռ:'C~������ٳɓ�,�Y�����?bi9����쫫w�D��e?�����Ȋ��k����x{�с�O4O�}�����&�\n;:b��aV����c#/|��&<�J�iW�
��E��nX��w���Y�{�:�Ǣ��d��3���������K��?xE�+n�z˄���p]JJ�=<<�}���I��@t]�}�(�	ƧN]��J���i��h� �-����9Jۅ,��T�D��w-��z�!*y�.����⦠�Y�A���75x�|zGf�}U�*�$
�f�jf��r������b����ܮ;�Rrr��$"�x��
�ڸ��c	f΃3jķC�b��n��4�:�o�Ϋ�!�<z3�Ջ��Y�W�y|BdD�w\���FC+%MC��9����j�|H�c� �.�]���k���|�2�Eέ�p��c�<���OvBH�O�2�޳g=�F�\����ؽ2����D(�
/�<����J��c��LՕ��&0J���d /��vR�����p��^%�YJm�K9�7Q6~"��b硺�P��]�kq�y��� &�:��1���>�s���D���\mE��k�I�ׯ�̣aqz`K���Rg^�nȕ�pq��XkZ�P�3���u������������?G������Tw��7�������uu�Y��;NM �_o	Oo^�+c�ș���w�^%&8���I�`F�r�t�����?$"�M�1��䜌j��Mٶǟ��v?�QN�V���.��`�!9�� �F���0���p*�!��Xb0
�z��k���|3���r�4���%��&X��������b޶��|i�y����V����O��-��a���l��Ȇ�ߞ����k���r�i/�nc=����O��n칁���!�%�.|\b�؇ �BԲ�'RO�a#��6 �Yk띃R
րc����^��
��}w��2��+�SUU�zy�J&!�y�ڣ�"�
��23kGpY��a�d��Sύ�����c���|R��]��"����QVz�l�V]�¢!���J��FLl����9Q=�y<yּ�� �2a~�yZ`����ϋ��KV"�}��$�I������_�ĕZ���b�9w���Za�7�H^	�R{E�tp{�`_���*�����UG ?�?Ux���Z����S&4��=���n�dW���r1�ަ�D���Ŷ|��IK�ù+-�*���<���ٯ�	�]f�ԡ,���jq��/���n\����!�tw�q]�	��^?S�r�qŵj��'ͩ�<;u|�D)C��۽���==V��p�p�� ���v��>_֘����8���Խ�k����Qn���R3ۜ�FЙ~�\\M&6Դ�RJ��	v�ڠ��3��n ��Y����23��N�nT��Q,�{�r��u�^75�
�$���Sy�l����g���3��ź�����6��m�W�����W޻W�n�I;w����H 0�a�Zi��ګ>eJ���+�1��C��qv�6�u��R®�eS]������_�-�RR����ZB��{�>p[�p��Դ�Z뤑O�F���ovw����7w�O������F����ּ��QR��r�*�<+��bF����?.�Bއ�\�2�E6�Z�W�� {�̰ צM_U���Yp��(�>���x�;���}��8����y4�ת���fF
KI��z:��Vޝ�&\�-�;�� �k �Y��uF�����h
� V*�޲=^W�!�;ʶ��n��gP�KȜ���b��6�6qӼ�<�N=���x߷o���{n�_%-_�\xƻ���ZU(U��'3bg��Naam0�77��Z��	%�@������\~T����tpF����h��L�>q%`ډJX�ރ� O���9��&r�S��̕��/�&K�nnSp��T2�-���E���C��	�oj�_ݡKE�S�4��$J��o���uFa϶�;��+������7��,đ������aaa��*�uaPr+�� ��D/][��)Ҹ��.`��;�P�����i�F�̃�*Ο��X������Z�	�	޸�=� �]/!�fb�W�Ac�t7_$���-�)���tחv�:u��wX L�a���[՘�����ҵ;D�Z�P먗)?��[!Lv��B���}o޼I�OI����"]�!���,]���3k����5;�ZՈ�;R.�ps�l�H��.��� {�ݼ�eݦ�-<�uWH
Ϭ���[R�D)@L@����[��v���G�IQ��[h��(�����5	zX�EK5���s[��N@y�ETRQw,��|��x��3G���!� ��WP������1w��c7��w>�M������bM�$�NI�d7�m�8 �s>��f�z�f���l��,�x�s� �,�+�G�j��1�欨����{Sjq	��G�����ul����*Iǎ+��ٳd,&M�Rn������a6J���%���bn&�8V��˃��n�������&>������T�|�ҟMש��EM���C������p��)��~�����W�N�h�uq��#/�CN9��J-|Z����������jC��L�\��.�;U��fA�}ܪe�<�wz0@=&�m��_i�M�/<���7�c�Wx��2��r��7&6���
E7qqaKRO���^ęW��b׶V���m/��3��ZP�=(Le��� %>>��*�� {����]Ԯ楶�HFM�dnW�����Oy$��C2=M����>(�pǟ������0�a���N��9�����fW������J�����aJ��,5īg�O������@�8\�Cv ��_�b()?L�|����Z�g'��ĭ�Fu�U���xԸ���P�h,����x�;n���m͗�����g�/h���nQU�����>u���4c��1dV^d?�(��Ay�o�`Zj`�E�_��~
g�[A�QG��#jH��T�����B����� ���o����yl6��U���fN�Yy�h?�N0�ڒӷ],�q�(��[FJ�����"��(���� �L��L�Tc'F��WIdn��:W�uq�q�Ë��5����w \N0HE�\�n��0�1�۫�~�J��Q&n�t�,^m{S{5��Ü���{�;��kjl��<�V�1����Q�wkv�ð��ō� J�l�2Xw���@�^=C��J�I�����a�Z����$��
R�c���#�FT=\�[�}{�����-ʪV�q�?I�@G]5���xj?������߾}�7)l笛��|3�w9�d�v��Y�~����S�MR
i�s1S	��uӍ�ڑJ\�}�QX�Hr^Vt&!oª���x-
ΦM�p�G�{��~zLh�`l"`=��lT�0��[#mb#'X�!�R:X����0����I^�����l����qxL�e4��!����>u]f��*�|}�����l4�Â��f*��%��QG��my�qe1&-E�������4��X����S�۶G�D�Bc|ܽ����<�	�tn�_��i�-��.��%�F�"����(�(P�H��-`6��z�>�-X_k������6�5����mUR�}Ѿ��5���2�1�R�k����l_zwb��*S�l��n98E�:��[q�G�r���d�N�K�4?9]|	�+ڳ���#vv,.�
tX�2�]�_fK�`Z䱎b�mYU ��������q�t�Z5@
��YY	�yh��7~KV��7L!N���}}��̫���5��c�gx�/
:y�#����/w��t�L___ﹷk���y�8�j�D��4��eْ��?S�t��IL4�b�Q=�����V�޷D"�\��N~�4���^��v�8���K�峗4u� �m��4dѪ+�����w�G{C�i�KYhP=(���7	4?���:88�Վ�[��0D�}w�g�ͣsFAª�^k9w�K���Bb�n�����ag�b��|.��Lw��f��"����z$�,�H�"�e3L9�IjG�}g'i�|���%�rPJ���|%�"��֠sq�s� c�R���j�􆑈w�s(u%�FECϫ����x�ll�H>U�u�������X��6�ڵ�ť���&Ψ7���{�5���J�O �ߔ�3N�<��&7Qw-�cu�c�!�$66��A3J!`�������;�_LӃ�I��X�n��$n@�;X�C%�_	A�>�Jm�9z�M|.��bpHȝ
�i��KnL�?"��n�c\%{,�<�FL�������LK5�e�f��
��sއ�6�AKrӑ�=fݺ�=���qwD�Hn��nl��g�Z���*�␼%�v�wf�~.�T�G�$����ۍ��+ށp��<���*�1�I�EKY{$�׽Q;�ck�����L��@,x�b�NI��[� ����5;��R�O�I\%%�ϪE���;�6�ߘ��dC�S����Q�S����!	:\��+��4p�<8�3jYT\
Gɹc$��JA5�'�O9y��\���4����֮��W޿_�N7�:C�HH2���vP�eߍG#<�]:�I4����/Y{O��U|�YWE�c�!�:W%-	,��v4{_�m�HSG'lI����Z�~ʫo�Q)-XY;���,H��5��On�uy����6
��N\9§�6.:��{�ܰ=�z
��ql)��vG�U�o�ɦ<��1ו�ڸ7��]�
r�߱5����g��~�(���㚬U��^P��~��>��+ <������������T��[FF"w�>I}(]�_:|Ƣ`�D>�,9�&�7Q? �4Ϻ�f���V�$\%LbpW
E���Z��@ܬm��9�*�͛7_g���ҵ����sߔvԕ"l |�V�fi����W�j��������.|D��s5���,a�_�"�n�rh��PL};g�7���st�����[���Ԉ��'cVkd�o�4 �;|f���M�i������ ��"��<ǝ<АR�S���֗�xh�n�	�>���l"v֣�6�����[d����D��.5��̘�޹�����$��HUy��Q������3�q݃9O8��kr�)���b��U��gʰ� ��Lm�_wh=EQ���:��Oƾ"��-�r�x����Q
�J~�9�މ��w��REbvS��/���^7�Ng���1=s��H�e퉧BY�]�z..��J Շ<V��#��_�U�����	�:J��Zp%pO��D��΢f�#Ik���D��Q�(m��㦭`��ٙ�]_��i�h��@
�U.G)hXJA�IGqt��f�I��>t 8ؐ�%\�2�1'��g���j�A��S�|'|�P[6Q�h�Z��V/]s+؆�X)���BMH�t�b�Q��L�Q���t\�gE�z\L���r�9�[N��L�?4
?�c"~:�UC�i������ooԅ�#�]�w4�_�O�O�;��b��T=5-�:5�$Y"W��r�f���j�(��'}v�B��t���찟T�fG#*�Uf���Ӳ���L||BDǱF�B���P�$&�~Dn���$����P������	����7���|�F��h��c�F�D��c��NAl>]�Q7�%�D�ϯ?˘�ף�pk�|��i��]�嘒M�&�uE�Eužg�Y/��A���ě��bbb�r���}hJC5hV"���b��sP��L���*n��w�Ϗ�^H�d�<)8�S�.��/Ɉ�Ӏv���Y��,�Uz�챌ª �y���P����_�?TA��d�dqWe��1�^Gg�������¯�w����~'�qtbg��1;g�oGh���\?66�BB�A�<q�'T�m�C)�s3)%"��<F\�Zm��)�����c>WC�O|
<����]�����,����t-�;���|_txKl�~�v�?{	L�i���ƾ��_~�Vf���� B�[���?�����y(�@˱F'[�J�}I���x�А:�n�ho�n7�VB��������TtNWw�Ӓ��>[!9�YG+�O��D�2N7d13�Q-ز��ԟ���s&�&E9��|�й������W�ª��L�Ѻ���:T�&���V�z����:g�$���5n�+�n~����^Qי�F�ꘓJc�5��OEP���֯���!�+_������HJ`�+�B�r�써h�%��8�襜�o���~����Q�=.:���LN����F�)?��T�P�h\�sa�# �$Y�n3jKc�GV�͈��n|f�v��i��T�T<���!����Ց�%�dbk�;��C���b�˰����0>��L1��ЖFc�j�vߑ �W6*�f�=�o�8�Z�u���*:,�ڻ���Xbl��R�{}���,Z�(�?((����l����qb�_K
�,��A5��ss(lE��,�B~XV�Nq�����!�Nޯ�ޚ�1��UOff�����L;��3S�Ae���)�ha	�4�n4�BTՋ�ꌣml���"7R!j�_��S���M���<M;m���:�ݤ#��v��AO=�辨��u%۫��Yy%�#A���y��k����nX����M�3K�F
�t��K���%ܺ_YZ��WK�:�b`��� ��y��c���P�J�LB5?M��Y-ۅ\j�!�?~�u�'��8�2��Q�]�t�W��s���BSJI�[��77�>L%{���57h�z�zR����7:C�m�/������}wͶHb>�1[wk�o�B|�wW����v���k�Ν:rM�J\mD�7{%�����0������a�)��R?z����M\_otH��N>!"�Ο����MW�d{���>G-��FG��"�q*
�^^rf����gI�o:XГ�[_Df��UmkPҨ�;qTG�c(�:�k���K������S�X���
�݋�!~�e �2ԝ��s�Ƒ�M�SG&Z���Z��%�g)�DƩp IΥ�@8�i{P���^��f#L=�:�R����W�Vw���pt�r�퇋bߴ&���8�s.9$y�N�ڵk__K�]����D���!ž7��F-^�;��z��E�X,) ����8��S阘9_��}2s��۾� T.M;kl������Q����7�h���KZ=.?�q�ϭ-C�:݃�{�4�!�d�g'.�I��Z׏�\���MzA�o����޵%�+K�A^��'Զ6�6<�8��u*��5�Q���OXqf�sDa:�1e��`����WF(�\����è=�������f>�4#3�y�:J��7O(Q?�x�2u�+�W��*�qUJN��~������Y���H�[R^��V�[��k�����@K�$q ���9K*0��:!���摒�r̎e�c�jqۓ��-�ܞ��r2��֮����N�e:�گ}�(��ǜ���Ҡ��M{Hh�ɾ8�l��WD:��.�j�Zb�H���(P�4cX:u�3����녜{����M9�����k�E	��ϟ^�����3!�a��({h��A0����ؑ�a/��k�b$<<|����(pzvx۠3kk��g^�2����?��tO�Մ�}P�\�r%|�M��SeR�Be�(���6߹���6Rާ�yVd,��p!�Cr�e�SS��G�^{�J>E�Ѯ0���N�ϲ<�a�Ϭ���
�T)�_[0^ w���*��=�*��:�x�#B�VG�V��g;Kp�<�;� Gm���h��k>�;Y=b���й�ZG���%��6�����?+T��<y1��'Ȥ��*��RH!,�����K�B�*:��u���6q�_��۩��|4�e[o\w������|J�Q�O�c�\l*�.	���B(<���An0-��Y2�@�~�Ź�vΎ���F��?���-+Bcj��������M�V����TQ����ME��(����7�~��]՛�w˹�cT�K'� ��ի��2�V�O [�˄�+��ߜ�o;pM����WF;����A$����ڃ/�|�P���\L��L�	yN�m<��S�'�e#P�����V�Ѥ.^W�9���㧰6��V��Jg�� ��ʧ�M#�7�����������mɱ��G�u����������+.3f����G���j!�g��v�����\�n�'��~c�n����y���!:� �&(%%�^T�����$�b}�٢F�Z665�t� ��w4�D�����H>�ٳg�o���������K:�yl.�������zF}����O��":�~J�җcU�雖/_�'a	�]@���?��C9�J)��}0���9Ǜ�O��{�TXZ�f�k
{�m?�V��lv�� ��w���{��P����5m��K=!���y������Y��3�:����R��󨓴~Fd��an��{Ҝ5�N���$�7>���������X#�����]KEݚJ b�=�r�SnvH�vӜo��Ȣn�SÇd���Ә�Zß�&ݮ�g�db�2��� ϳ��:�@��R��y�&ř�(�9#�zO�2ݜ����ݜ�(ތXG�}�rS��a+��*�����Cz[�=f��V�	�Jڳ�~�YA¥]��VV���w��5���J�Z��xg�Q|�i��T���H���턽�aR�T�����7OeDV><E�6�}���S(�`�2τS�@�mE�ij�3��a�|�:$ں#�)`���q.�n
�ڻ�c#�4d=��7BC�5��xWϚeBt�2�vj�T��ʽ��s�.6G�U)�3�Q ��b"v��Ň�G�:='�Ջ����%�	��M�Q�s��B�OW�~�Z橣��� u+I;
���X��V��>%o�;��ڒv��L���.6�P(D�ӧ{;�'�������GG�X�W��>��;9z��� �7���gǌ�v\9��K�LL����+H�i��o�QJ�kYv�;��iO�w�'��A� oI�ۗ3n��e����:7Z(:D�Ŭ��W޳g}��c �Ҍpt��@���3ڐ���s|�,�:ِ��/7�����W
�}��E	?�,�C�bBw/H�� ˺�J�G�^!�z/�Txz�F<����#]`ް���0�Y�d��$iiiGB)RqH�nx�^�Jr��<��gΞ�@͊����
ɟ�/���w,9;��ҧk�l��;w�urr��ۈ�3��dq���g������uUp6Y�|ty�R�����gf�<5?(��ky6�����uhֿ��^QQa	�s��0����H���9�"�b����%ps���Cg�}G�@!����0<���lgϟ�7L/�)+/?؆����L�uD�
r�p���>���^()l���F��d
��<�7�~�X��y��|��yk����\HO!�u򎍍���u:VLL���J�J$n=5�}��Av-�ꮸ9����и�nF����5��������.쨾����TAv�T�4���W�o�w��.5�j��s���~%i݂$�� �΂Q��p���0$�PSG�^g�!��$���pmoEZK���.�g�m��m�6fm�Bz��7>�~��Q���@�% ��_�=����[N�����2^�V�v��SUU��<���A�)Z7�B�V�@�̶|Y��#��T)�6é	��� �)Aļ��^����(�ηm[0�N�_B��̘Vz��o������Ԃ�W�k%~�GL��@��H��a����������`DRRR�YFEy�?�	.ɗ�փ�������jN�(��˗R��on��-�YV�A���ו{N�zI���yѬ���ԡ˂:\��u������B�qTҟ�.����Q1�Qp��H4U1�`brGZPm긁YܔơCg���T���� �I��_6oJc�)!�kV'�6^�E��#��6�+��&�_�(� _B�\Zn�� �(�`���}j�K�G���U��*b����:��>8���sq��M���@���uJ��t���c,~�С�y����*2��-��{���w�NK�BI����l���p��BQ�xO&a����%#����;�v7w��%u�%�YZ�ݸ��&��M+�Z^^~�Q��R�t��[�Q�n~�P�~�p9���P�=�1�"�sxP�ߢ��m�j1̮���̶\YΝ�z-�:&1��XL� �{�\\9���S�~y[�(5pi熩8��&���44��� fjV16���A�,��?��a��<<!_�|I�h���b0�A�����kj�w�}ā���}�l'�b�`��Ԝ�qn�vC]� �9@�9c�-�gp�߹y��%�zzڧ� ���VЙ_��읰+��ۏ�m?6���B�@)��(Y�بӏZ����%^XA�_H�v���۽��V'�W�Ӆ���&��^Fٹ
eeeG��T)�RZFٴj��ү��B/� ��UN&q��A:�-��B]�1>�t�/,]Z�c���i�
][���+�Q�,,g�n�Sn��d���t^���W���#�2i�7R3G��=R����/`�EaeS��di+R��Ϛb9�w��4p^6��P���r�C�h݋��J��2���&ͧ)~Xͅ�@�<2=vb^����`��v:9pbn���&-0�LS�n�߿� E�Bw�];i�R��}�d��cSN���s�^}%Fl�6��4�Loȧ���8
�d�w~?l{a�L<��y�ȭ )i�r��~}�4�A��+{>En�$�8Hy��uZ�⯒9%@3��.5�Ш��f�+��B�'��E�Y��T��+���ʒ���}��;hSΨv����r�ԫ��; 2��9��:��F�M�]K$9ڦ�͗Q���+�^��+�
� ��A��4i,mk�����;_!����2���0d���Т��`C>W4xߪ����}'M��C��p<����Q]�5�c�`yB�[��q쿖gDWn^]�w��(?��n����0B��<���!�cU5z��d��ˠ�j�U���y
�י����y\o�pD&��,�U�F�ϦG4�>�Zp��Џ?n޲�}ѝ���W1F����B�������r���$�j3�@+ێ���\4����y,m����ķ.���{TYL.˼
0�¢G�_np-����������w�jYAB�F_��� �_AK���!�CV�����;��v��2�A����p��mXOs�U�N�ظ0��Y�D�D�߅/�)�9�P2�����Ɔ^�z5McQ�{��]B�� �XX���C���y�`(HWv9�'6/:����#�1����"���ѡB�[n?��K������p�e����t6��|����Lm�t�A��v��ST:�4B�翔������/9ܞ����b�RÜ,���ѿ���t9��᷻G,�n��'�.K?��jҹ�8.�xu��~�yA���vs.��+My<�B.�7�N�z���v���Ͳ��Kt�C;�i����sj���U�Qbtg�t:���j��)��Vq�KD�]�]:OD�nĴy����5=eb�?zb�◜�c�G�T士�=���k%֞ke<_���$���"���.�������.��2�~1ap�e���'Ht]Ѭҿ�O1����P�)f���EzZ�T�����T��������8�U�
Lmd/V?E�K�@b�����	f\�0���r�JX��ѯ!�:�j���0��.�q�2�~F�=0#&����0÷	�X.����U�3�3,2�q�u�=��x���K� ��W�nlg���3
3*1.2��3�ѳ'S���f���k�Z(r�"1�ta ���|UV�v)��%��s�>�*�,���\��bA�(��ۆf\v�\/,��e�}/��9c�b���_5��j!��Sn�C�V���2z-i�=�/���z�g��u�/+�}K�r���V��8��7]����g�/<cgx���]�'��`�f^7����b否�0s���˚ˊg�69#�����b�/���Z{��Jѿ��R1S貢�]-\&�m]K*�`<m���`��,aM�r/�O�?/x��ӿ|����-�l}h1Z.�ni�S���W��n�7�d�p�%}B9	K�cg���3Vxvօـa\?�D}�癋2�0kf�aMa�x�]V̔�k��6w�Ҿ���K���.֡t�en�Z���I�h��&�� $?���<�ѵm��|�6ʠ�R���-m~/���IK�.���3�g}ց���ZE�����=�o[,]ћ��܋|������_�����K�m�T,s]����L�C����t��r5]�G�;���q<�q�;`�^p�l�������f�J-�Qۇ.������Ӆ_�yI���K��[��k��,� y,w�J2�)�R��M*�/��`�.;�K|1��sY�,���=2�l�Z�'�Le�`B*L(��>a��sS��3t}�A���g;��΃���m�����4(��tY\ALcc�g�703��d�}�Ś�,,,����� ������PUT��?�����P�\��1�|����O�09�����.����g5V��d�i�Z�OB��-����-����-����-����W,ɲ��Y�����z�O��w��{�1��~�
�ʖo�?f#���[�o�����Z��S���� ��������-����-����?�#&�+�F��+����´�X��Z&��/x.5�?��V!��q'�c+��Ά�o�11[,Y���
�n*�h,T	��{$|��U���ޱ��z��|�.ےDl��?���rN&��ҘJ��l��D.��6+��	j�В$/��sd�%��7��23��;�"�c
���ma1+�w���q,/Y)�2��\ϸ����1nc�
F�\�_���"��-��E䕀'�Le�����L��-�ҋG߉��e�ϑ����������Ϗ=����XǓl�_��D؊������"��-��h�{�/�x�[���̲BEWWל{��at�97�Ѱ��H�ɯA�����~~O͐xt�c���<g�g�nnv'��B�ց��::�R������^_��ᝣl��{6�+�̵���T,�pW,��'��u��*��c9�(��0Lev/Y[�lV�"�saz�~hc�� k�4�5L��jd���0��d-
c��=6�6�+���y;��n͊��_O͞�������{{^����,ӫ�5�x��;�u�Yg��;���K����-+'�J�R�!!!'�1|�@o��[JpX�rrȩ��������MJy�݄��Y�ߍ����!��������q�0>_�w%n=�Xq	�Y�p�\l(��]3�D��JN�n�5/�OOK{dZ�1�7���#?ÃJvdTZ�Bں�A1�Y�7�v��K�FW��}���������Ƨm>�D��k�{`�ɮ���"n�Z�QeFZ����]j����ڰI���8g����I=pܽ�ݝ<�lp�h$�l�/՝�zIN����*����F*�>�aɼZM��V����y�!T��,WN���oq��da{�����5.�俬�ɞ�a.��"�O�(��(x�x��M��ZP�������>����Y�_�o���-j�C���2�����ﳖ$�Ą�c�]�,mqg]]�x�0'��_���%arx_�]>��Ŝ�Q�7V�jht���h����Um�3NC�� 	�LU��_��^�i������X�e��LL�����0�h���Di�,���.|���3���ljb����N���𣲈IH$=�Kj4�j3.�Ū����a�g�0���t�L9�kI���N]!��j[è�9W�#��1������Z]�/o۫�g�3�����,YZ5�̞�8sé��~f�1ƺ��Ə���<����B��v`zr���uC>�v�%����FJ��vf`X��]�1�[����{��^
�1��ˌ+.�\���e�aO��"ɐ%J�±�L��
�>A����]���;��/�EEE��J �VHBT)"VzQA@���  M��@("  MB�TM�$A����>�+���;�ޛ�3�{����g��Z�U��>��c�,lf�ど�{�q8WN�F����פ��Q���5�!qK:<��Q��>df��S{����n}�s|Q,<hN���\|ζ��5�ϊ�6y�H��n��C�̌��I����!�D��O�ڼNs���u��|qN1}T� Z8~�ڀ�ps�d_�E�}ƭ�9�L�(MAt?�m������OK���R��̮;�#�x���X5f\�9�b�v���u�r��h/�Hu"�v�`���۟�eqK;_��Ґ�	�+~�U�
5��z����Uz�-;eh�	***3�l2q'fW�"Z��\W�{�e �d�&Ց�C�544��h�;��dK�^����a������#���l������X�?���Q{�4ొ۷l�-��&�j\��D�hFn�WNf��؋W�I%Kv a��Y5e�++ǚ����^n�������ʀ�p$��r��ax�H*�����6�$����𙛛;..~m����c�����&��1�b �b��aaa�Q���щ�0'�e�#����
��V�=���S��ƅ.�8��H��2Z��PiJ�fQ`x��YjJ��!�����.��uh�Z��f:�wB_��)�c����,�.-̨��8�wnrӯ� Wjcc�\'��'I�	`R�J�:L�o����G�c;���ׯ��6ˉC��;���Ϟ9��|���lh�)�0��Z�;up�ɭ[��yV��ENM�0��{v�ݽ}[��=.-�c�	��Tmee%�N�����Ǭ�v�[q�4��l�ʝ��i�6��R�]�Y�[лG�"��J��fY��I
y2����!�ڵ��P�c�Q�h ��*�M"�n��&�� %���q�����M4����Q'��jMl�$7n���?ݒ�s3Y?:��:S!|&��\&����\]�Ki"���G�>~Tl�2�����엶]9FtĬ���F2�및�,�A���c�qPK���� |��%�fP����Sf���zNHC�M,Ź;1娇g,j��@h؏&�ӻ,��\�[��S�A�� ,S�>p-�6'��DI>w*�i�6� z��b�Z+�=?�NEQ@8 '<G@~�l�!}͹K�$��J�����]�(�����pK�6¾���\g����/1���Du8�#`X�]b �,�
lF;����6�Nc��ܯ�>�_*�A&A���p4���{@3���<C�kNP��>�mH�Ѣ�/�K�ǆפP�rm��6�XYY~���??�r~�UF;�f��3�ʦ��	�-<C�e�U2�kenJ������)����)�<
<�sD�a���fԮ ���������c� ,�ꕑ��q���ss��0]��� �/�45JV�g@J�Yc�v��ӫ�R8�3��ƻ���pE�~!ʠ���~(�{2�Z�*̥�NV����1l���M��)��]�r࢝Z��R��N&���q_sw��S��7o.Q:6�6�Ji7X)퐡����'�切�4�S�)�@OHH�B$j�GF�v��/@n��"��ju�.��%���@8ӥc�D���;��U��<�z��8"����L-,ِ�y6��g`of*[��|�� ė����Z������GK�����d�}ޤ�"ڊ`c���J���GK��^�n����aO���Q��ٚ� ~��nC�P���:��q���U��=h����&'l .7��&���L��K,��a0A#A�v�Omg�'A�qUʛ�)'k�F�� ��{���E��p�)E�"CK��&�P����*lԤ�~�2���@�Sz��Q�k�;�U�@K�j�8VG΃��r��s���E0r�v`��7O���\��ꚲ�di7�?Pʁ��`���O�*\6�*����e2�x�c&
��Y� ����*����L�1�iH@�S:_��:Ps�$+8j�����J��穧��8�l����M�Y>�2Y�p�ٹp���#��-:�@E����wg��~E����#a��m/n����O/�x��9Y�ʳb_le�Ϥ,�u���;\�x��ozU�[���������7���}+��̘����@��TuW�;\EUu���kRz�|��kN�q���F�|t�;�?Z��Y'
�/r1=3�mc�4<�S5U-މ�-Y��\�lP�N/i��#,,|�J�۷k7�f?5$��%�.���/N�O���F[@5$�����#��]��������::i�\�����:��` ��Z���/E�L�H}=�(�����.+H����)��9��~^�y���R�J�爍oi�U��;Oꤼc~V/�z������-6��z��i6��[�̞���:$O�J�ԣ#����0 �+D�ΡP��!)�uDb�X�Ɂ�س���M�ɫ�Z�����9kamt�%�n�_w\we-��g��W�k�x^nƍ��/g���Z�oU��^���Z��]�С~Z���}l��^��̅+ʭ*� J�QTvRP	~���m�~8�=[FQ(�T�S�f����R��ii�7�&�;�ٮ�\w��=���p�	�q΅�����6�gm��/7��eAh}��0���g*�F��eh�D9�AC[�.f�q����X�^�����g��<Zj.`Fげ��.�8��:G�a,f>�������%t���(e$��^��_:/o��T󯫻\��qK9].((��()l��Ɗ;F+g���,��	fH�'!���oR�����	Q���`8�+�v�3�C���l�[�({�����R��m�C�HZ�ڮW/żN:�-���� ��Ҋ�cO�x�GGF�޽� ..��/tUQQ1"GI��_�nw	')��n��CE��w4<��Ś���d��6DM�����4M��qo?�Ab}����"nd��#�n�sFR���QR��i�-r�-�ho�]���3�V\���SA3�9f\�n��ɏ���LMB��v�]�v�.�k��9}�n:�]5r3���N��^���I���������c�^�f
@u�4�l��G��_��Ĝ�%����]jg�G��'���\����YŒ#��:�'�9��B�vx���T���be�9R��ho���B+C;?ڛ
�ĳ�z����[ho^�NZe��+�]?��<�ia�Ww�-�u�&��o.�Fd 恜>�˙�b���p��̼�1��a\�������6������\`X!@����?���ڽ������mQߞ�b����<G�;=P��7k��,���h���"?�����~���CL0wYr6Y �6��w#�`��D?�!���m��oۢ�u��7q���������jjn���ၽ:��F�.]�����m�;[j��CM�{]�z�QZ�Z>G�5���#x�a�mz
�t�,�,�F]�gF·�I�݃��(���&V�&.� �-�������j�mx������g�ڈ��SSS9�T���4�;���[^�	���Hr	,]	�6A3�/�5���۲礧�6}�r�`M%*�lOy��>���F�[X�8��-��1��"UUU����)v,_���|g��t����"����eM������JB �	j��k2��FK��a2 ���)3+ĸ�8��	_�R̊ۄ����l+�1pp�:{`ic��ֶ3�l�:8��޺��@p"=Pu(P�@6��},�H̷M7Ebs�~�Yy+���* �?�~�������A�JZ�����@�Z�y{r@@ P�V�0�{�?+t����-Е+W����
41Lvn����# Ъ�m�e��60���w���i###mi��a8h	���p��b�:�]�5aC�R��E��Î�� lF���@�.7S�^�n��������$��U��w�`�4���8bz��Z�y�1W�R;���g�-�9�� H���IT'W������S�uc����q�!�������"�3�pX�<
l��9��d���\)M��
�&-5y�5��ɏ����R��>�!�T���X�X�?�w;Z↾��#��P���<�;�����k�.�V�G��2x���7�����H^��F{��J0�܇T�\�s,�̎Kq��3�6�~�FFR�5H��@�LWW+�����\����[{�\м9Ͻ9�s�*@�}wPՉ�J:K���"9X�:5=��f�L&D��v��e:��)Q�O�:ů�>�	��%�K���/�_¿�	���L8_|@��Y�����K#\��Yz[�<ǽ,��?�����O�=b��s�{{�^����C������=�8�pr�{�շYR�e�^�8�SMF��i��6�l��{eA5��<iA�T�e���>x�s�Hy��㿃��z~s-Yi	�Yvx��&�j���!��m�O׹�I'C�����hF�ű���7�l��8m׻(Iǟ�%�M��c�u����s��3��^�+�j���w��v.O��|^Y(��X�t��,U�	�(ɹ����^?����ɁzlGj�+in���~)6��[����H@��v�	J�Z�ꌢ�/�"��%*�n1}Lϋ߮$j>	@m�\BV�%-a��V"�,�����qn6�8�!��G�fZ�h�%��}F�8���/To��By�!Ӌ	OJ�+�7�<�8�N/D�m�#���;]:��+�Ul��*���Yp�Q��;��SW�1�q�-Z��(RaǪ-\'ܖg�d��w�N�m���Lō���L6���p�Ί�Pu��Jq�\�p�E��w��D�-M@���j�u[Y�7����d�Q �Yj�i�~.,����]s�l9�~��dȠ����oP�4�f�'�f����������\�B���n�4 X����uW]����>��[ˇ߸)
���U��\��V��)>Jp��IoN���s�n��߄%>�X"9!(��MKU�Z��sB�N{��d��Z�B2���I�)�nuu�8��B�Kv�${�	I�e���(�7�wO�5��b"�%'Q]�h��w�����Y٘"ϑ9:�����ֽ�K�\.��c�Itpc�J��般𳆲ҥ�?��(Κ#K���pF������ |��3*�>CG�O.��9���"Y���E(j�f�3�~t��������(}�=Q�4��t4����!�8���g�;|ź[����8{��t�E�sf�����}�����P
g�Gm�������<�ʂ��X�	-�Di���[kRh���udK�Dѣ�p��
���Q�സ���At�\@I��7nb\e�\kM6-������f�mԤB��Hw#:B��Ɉ�&+����+sN�C<�h&6R�$�ၾ����orD�LX�u���1t$�	g}��t�k*Qfi�f$�����4�_^���Gut����}�x��s�'�w^��j�t���\��̓Ϋ�%+�΃t�v8�^�Z��[j�r�����~#/'��,
J���N��!�����/t$EI���q;�<��[����H>�����/Y�<+�U>>��~i���+�TL��X�����d�9��Ɔ����$n��G���L8�dHr�M�;�l��b.����P��7Gad6�TJ�?���Q�����c._(�PB��3Ƣ�ua�a���kD�1(��'��z�����l�]\�4�5���;���#�#//_��T`��aNd�Hʙ#n�e��c����OʦϾ�r��	���]�,{��� �J���')�
���s� ӻ��_7�n|*DV*۳?����]�k��+�&�! rM���$��@�W���Rh�O�݉?��
x5z�қ��(�`Ei����?&���T�P�D!�rđ����N�{��4���ch��<Ԁ����*U�珡� ���&Et�"�D0+��#Az�ط��%pA���)�?��]*�#����Y�}t�t��協B����A���o�AR�Q:M`�鞣\��y9�.W�ߖK$/�_����Qw��yxD���c��s���Ӕl�e�,R��	Q��- i���&���6�Ku]�7���4y�$_J�dw�B2�H{`(���G֓ ��K)tȪh��8���H����8#��� lXȅ�%�6�7���o#�WG@W��m�gu�mAJ��XVG��QQ��:�(���l����Y�G[HP���y���,8{OJ��H�6�2S�ML�K���^ʵ�OAk�I��갤��m0�
}�E2ӐM��SK��E!�H^�(��f�}�j�P|Q?��{y��]*��j���&�4�!x�/�E�w�%�"�
��.���U��h��l���P�-2<���$�oNUK�_T-1���Ѳ"��%V�/%r.�d�<@���ƽ�	�IX"5I+����5r���x�6BVU�	��\�I�&	P&�:v���H�yJBV�n��Ra�:~U�f\�o���k����!�=$��-�}A���/<��R -�Ց @C9B|�:��^��z�����*�_;0��mp�*U��Uu��q&�ʺ���KG���N��j��R�lR@ ���A4�4(2��� :��¯ݧY 	Q�]*�)��?
#�XJ}>�z��Y@�	�]Pu�o �=��ʯ �eZ��dQ<w�y�n`����A�k���	�hy��d��Ҩ[�����J��y�h�As)��L�$aClHT��~ع�'^j���*�]9�@謤�q�z�:�<T�S���3��~�IG�%�Y�6��{8l�U&��lC���:�fJ���)W�ZGg,���U�>�[��~K���yZ[	y����xD�/'�$����9��p�b3�_o�6<���u����Y"�B��
�~��Bc��
�"Z�!4����3~r���ʐ�����c����^Ū�tV�9׬?"�at��� ӧ�jgٷ#3\�s�J�nX�,��f�K���(���4��p*
�j�ي 9NMB3�ٛ�=��ܮ ��SU��{W�2����%�9䁒t8%�'N��[�_?Ȟ�%bx��/J�P1z��< Uxm�Z�����X���_LdE�Ʃ�n~V};/�nO��{ �5���B���r	'�,%��k���8Tr���pe�i�󼒓�5*l�K�<�3kG!ϙ��,��N���9gn[�*�\����u?8�+��H��L쓔S��sj�#��i��Pf�y�d����uh��҆[��D���Uc{=G.�y������Lv4�^p���_���-�Od��.�T����6��s��a��{ف������vڑ*��^�e�ʠ�Θ�up���hR��b��U=Duc�o�񈭼6���[��ߤ�R�o���t���W���+���b;7P#�,�j�ky���A�/j-i�_n�5������`���ʎ���	w~�,����[;&�O�ͭ�h	��7������F�m���\��dgΑϥ#ƞ�$[n����]�'�ʐ��%b&���|�"1[�1�ve��o��n�dL�V���������<���n�"�/���Λ��ya��q��r�)�R:Bl'Pz��=���w�]�2U%��g)�{tZ�͓:l���nO\���a�Ϸ���{A�r�#�� ���V1�`�UЌ&J��A
�˕+&�mv-,I��[��nܾ��;�Sa����(9���dU�G8���pl�E���$�����{����Y_.f4" %r��O�� �C����}�;��F���s6�C�Y�'���Tl�p+�I�����1�����g3u��"z��Ny���i�%��|�.�Ew���h	�L�M�|6������~�׌&�|C!���?�W>��C曟��U��5[�S�x�5gS� �FDȦ��BE�S�&0�%��=D�ﾞf����C�I�"��;J���;�DTU�X������3�=��:�����=GdU6�w�x�N����9wV�o�y�4i*5���b���Q}�E��܌��
]�t�@���UĿ�o�- d��4O��g�#U�>��|�v1۩I�V`���������*��>ݢ�.#Z���/���@�꿚�]��� ��Nnf��>�d�q
~ ��_�J��s<b"���z�J�7	��P�Oأ��:uχ�y(h3���n�og��p�=�����Ǌ	�4�-��)�jfʟ)��+�
��7�lô���c�_}�^��g2�7��d{�گ^���j�3�����g��(�_9�%�-q|�JPM*���8�戝%k����~�%�4 �$0� },��h��Y�şOK�;�H��N���m��eXs1E�*��>`29P7[)^�~z�b�p"W�&�	�i�`�7� cw �l{vL<,D���w��'�'�o�����@hېjc�@��F�ʥv���M���ǘ�Eop��lc�,9EKܠ�a��?�5OM�J��Tj��{�vU`IX�{�i�L+ã@<�+
6�.�8	Vd\�i��ԥ��h˺�o#2�2�K(l����	���,ˠf��,g��^�����R�����T.Z��G�����p�sߧw�ݡ�|t��
C.57L�Q�߇�9���#��D�_[�n��	1o�e\�/s˸�� ��23��	l��F�b�Ri���k�e>���j����6?��C�>�����_¿�	��%�K���/�_���	�7Q���Ф
��x���Y��Ǔr�ْc1�n+�SlkD�����e���7٫s���I�����jM�_�}D#�?:KNiJ��x��qv��h�����țO������a���,���_2���m:" ���%�Z1M�;�"�͇���F�D3�Y_��3ȦӁ���gi��Mu�`��E�U��hh*��ԁ���bܦ�H�/pb0|�T��dջמ\ng��Ùsݽ��������Pl�(V��v���u��}�6y��0ف�a�ӯ�r�>���R��$���^���XN �28 N~�8�C�/��T�k��Q *�(�5�Z��BHc���P��u@������͖��^�`�V �%�� H3�=�۷���[u�����A+����-v���|����/�ȭIx���0C�+�x���uz�������:�c@�Va�Hs}��74��!�>q �J&�V�V�+��o\���>�"�Q���7��"��5Qb���
��]�k�S-�$�����d��Z�k��;����1`�e������.�W��c�Z�ti �Y�5��"@,�m�����Za����jʕ�}T�! 7��P�%544��&�B	���:i\$ o_�k`��g���s��uՐ�V4z��ݙ5�F�uK���u���� 8�ϭ�m� k�����˿`��x��������5$P(ּM�}`�u�4V�~@ɿgMF^/ M	���}�ݏ�E��r�\g��,\����\f�0`"�.� dJ��7��c#TL�UR������%;
��=�{���D�2 ��)v<F�q �lYwp�E0���j]�g�3Q�X���g�>N>[�*@��G�$�{��ׯ7$$%���;�U[���l���7@�ZO�z? 8eBh��u��\Z@.n�5���D4�5�C�Wa�O�ɒ`�HE#���T$+ p� �+��q��p,Z�5ܫ6Nu10%4k\M	]ӛJl=�. ��C{�=���CO?Y��X� ���]��P��`x��G�D ��-�i�ϭ�� $ǁ�w�7P�gL���"O�C.�,4;�Q]�|��a^g���*�w�z3qîgJB���0F�Qk�J�}��N�H���o��?���د!=(t騴J�a���-�%�K��lE"��}N��a|��qMg��P|\���Z��ޑМ��[;"nd�3���M�����O�������s�Q��B��
��Q<���Rɿ�2���/ÿ��1��?B�^�ߘgH@/ؒ����[k{;V�<� U����z?��H��v�LNMM�,#2�h�U^��7b��ƙʐ����_�0,������ʲtrBb�@�-��xxj�� ���@�n^I	OKK˪C�=����� ��~�3)�,T��_\��?I߿�3���
v�JJJ���佪�-##���d��R'��!7*:����������Ia�M�R�(�K�)=H�����f��5�~�&��K>�]hl��֒D�˂�4=��3EhA|��`û�������;�s3$����,*<'����D��2����3��h�TUU��XsMEE./�T���b�����-�,��O�>YZY�T��8���եŢ{6�|�<[#���ttt��x�����~��4�-�<�����0���/��ug#�PO&_��_I�I.0r��r������X��veFt�ѣ�g��#���ܘ/��%��\U�xv��	��u�s��7vw^~�q��89�&�%�l���o;e�U5�97�=?D�HNLI[XyK�.�ƽ{p��zW-,�B����#V���Θn+\����ēG��ƿZ.�-7�B��}k��6u��;Yc�
����I���gE�ܠ1p9��ƙʇr�3�wA�����Lk�Fcn��Y��=��;8hu[7h��A���Ǯ�x�<�PEA[z��ֆ�^rCl̽�$��,<�jh D �N�Q�u%%��ѱCYn�	/����
dC"_\?������F�������?��^H7%+�Xp:$e���{NS�c�	����̾�+�]����^3�p�����1'� �HL���
������;,zxtFIA�Gq+~r�"�p+�;W&	&��*4;�E����ݬ-����Zj��-n'l�}|p3�n��[�z�|:�Te���iv�	���0�Ӝ0�<)m"��#���gj�IT�*���ɉ����s�sN|��h�ąh
j��D&�"�+H�F|��&_�����sDr��g<�]v���IH(�{��"}w���qN��A���"�W\N⊷�0�nj�((xq�G`��������{ˎ��d�w-��x���m+]	ߓ��́�A\�$� '"h�a��LQg7�/���%i���!���j��xe����[��}��+έ,�um4�>)�d��m`�p�le�����J��d����L?'U#�D������\�D�V�{{�o/���*�:ݹ�t�cՇ���I�!$�?r�W�T��G*#�d]�ud}&.��#��ׇUf�!;�_%J�IAD��;L�W�C$0)�@���])q��&�+�BP��aC3����]�$�?m�+OGr�V�|(��y���_X��mq�KO>��5[� 7��[
��o�zJ{�׋�������J�a�U����nC���4�Oq���*6���.��Ы�H���~��I�I��*U�3�N��2����BE%�ӑA���~a�/�h�<�y+�����!pz��ܯ�/oٴ���g��qI�)q���3o��꼹�и����V�9�̅7�D�%�I�<1W �8L���f�nD�-��Uyɩwp�͏�\H;��������O�M�����_\bk{c�*f��՞7eU�]���7y����c�Q�u��x�
�w��q��ȍ]"%��VjJ�s���v+�Z��F��A�a �(��t���B�.23O�OU4==�g*���	(� 1@�Fn�ݘ��M���t��w��Ê���C��^��K��g��k�Vxz���5]fBZ�dB����ځ��f�����;�{>X)�^s�|}���m����?q?�ī]��㨅vHk�O��K��~����z�����,��Xlf�?É�)�]g����'a����3��֬޶���3�s8����R����Bσ�*_L(�AQ_E63�6�=}��
�R�ZjB�+�MRvGøQ;��+������M���qwk����v=ͭ��C{e�/%U�Tul��7g�i{K�m��6�a�����ܾO͉�.a���6W�[V�����{#`z���&

C�T�//%��a1��	#�Ǐ�#kTwF?��ִ+o;��~�w�_Sw��G�6�*�V��)��o�MvD��M���֎�D�L��>��ʻ��s��?.���w4fRմEm��I���i��������L��M��۔ǿ_+�n9$b��,¡Ӛ�\�DB��d��H[��r}bO��Xe8��Z��kl�Y�s~���ȩp(-���o�������<״s�B�Rxi��N/pȭO�;8[~H1Ǳ��j��T�i_i����~Z1�'���CH�ś��?@!1������%���_����5LY�=Ly�ț����[ށ��Z� @��
y�{Ə���F�Y%��w�:��z\�«���l�y�?��j��sw�9D�f	�l�c�8�/�R�++8DT�.�X�\��T�\N����Dɗ/UIi74X��l�/49)��t]�*���M�z�ۓ⎗�ؒ��>t������~O*"|��e���od��u`�؆<����G�q�oN�?���#��knS���`^<km__��).iף����E��<E����3!pc62��͏�q����JG�8��X��avN�ZEv�L�|:������@�1�{��B��`��F�]��u��_�r�����و�\z�ԝP��e*~�e�f�������⤠l��>W�ۙBkS�񽐔BIH���\�)Qc9���,�w��"�[g�� }5Oi��R3.�**����H��P}�|�L#v'�쯺��8��N�r9[�X}��۷���V�I��TK���A�P�T�I��&ܭ�f\7��첩�0{T4��HBJ���}�Ӥ�����Ge��~�b��~kʭX�j��� ����x�9�m!Ŕ�J N�N�d1N8* 2R>�v�#Mw�a穂���+� ���w.,88���D���je���w�.X-i�<�e17}�;����/��pnyQ�k�ȧ���8�ږQ�M
��Pp��%w�ƆO�]%�գU��b՞@�pq(��ߣ>�Q�]�6���n�L��jG��4u �`�Q�]=�j�dd��i�K��o����\�K�W���%6���iRR��9G'd�T�xyx���wy�pb��)�Zsb8��6������Q�p|!�jRR��6o��t��k����dk H�$�ʳ�R��W�7}�?����� q�c@���l<��5���T���֢î�n<E� QY�߷:,V�r�`�\N��W��4#����"Y�>�*,Ǽ|pwG�����#���^��a���V��]3�|�N��ַ��C{�4>�%X�p
�`O�|	ʗn��c�E�4*�o�i)���Ywk]�Uƪ�N�#[��+�٩i7�޾b���������M��|	�wU�6W�-�T+l&ʲ*�~��(E�2��U��P�h�̌�l+0�����N׽a�`���QI�m;T=�NZ!-Mˋ"�#?I��_w�-�64	�|���ۿ� ����HpJO>sI���Fuff�Y�A)���K��]�'��$f� a�x|�T^��ԉK�(Y,��װ�Xk�\~�p�6jD}���]�l�R�~tm׀�ٟ3!�h����b�bN��yt�����m���ح�=$d��x�����y�'$��%YX�w�+V0лyЖ-f{$'���*��h���;�~l�Н�,�a5���'�5�Z�]L�����/"��y�L�5�g'�jK��dv%*�UWx>��?� /��#Y'@K���YV/.����а�u<8܇}��_�΋7��c�_h��F����iE
��1�ͯN2�������a���I$`��}#[�nT&y����\�����s+3�z��_`�BО�?�b7���#���Ğ�N�㕕>`]@E�WMSA@��{r��r�~rk������m�So�ć3�D���8���U�r��J.^n4�~:��,����Ao�r���2 i��P��G*�&]$V#���q��IǏ& +d�אoJ�ӯ���T�"�g��Ñ�i�@�uhܳAoZ%
�`�)��'@g�Z�D��_��	�a|�D�]Kμ*�Qԝ��6�~0c�8�fƒm-���3B.>�;���y�wl;["g�SI�ma�-�6�-O�\��v��(�\	.�(de����Qs��{�Ev2���(<��<h��M���ٓ�L �&_VA@'ƍ��!�>�?0p� �R~�5۶�1RoL�#�w*#���z��_�B�#� �Hjm ���,�Rۯ�Z���0����c��>s$����)�׈�?��@�v4�,a5�}���#N�H�G��8���WV���u�6���������ؓ�_3��<�Kj��<'7��l�5[��`�q 7���c����&և�32TTG��nx�s҆�2�nN@`@�H2|�:�<>te�R��f�y�.?,p0�S4�\A�	v �n'+ې����"�vݹ�L:��.o�H2�����T�����j������Xr��-G@�CE�p�+���&���&�sj�}��r�:��{���h�N��.H��U�������Wc����S����D�����zc�R,ù�Vc?ը�;
f���P�}mT�rK�\�a��7�=�k�ݯ��eq��̶'����=��#�0�2�3�ם~���sp�z����$��t��.u���݃'R���^��0Tq�����L���go��ƶjhb��	n{Y����Ր��M�MON�h������綐����&�P� �x��lM�O!y������5׏ ��e�o�1�ĄKUώّP�U*Q��7�]�V��q	��r#�\�`g��-=ofb�y`�`�s��;����
Vb�iK�y��`���Ԧ�J�5�-����J\a�ڍu�C;(����~p��a�t!�����e9� �u��V�P�{��p��ǝ��-�1zH�|,׺��I['[��Ĝ�ga���ϔ xGĸ�0�/��z��n��!#7s��ԁЧ8;w���Jd!�F����1���|S��%���'�*�'�����۴�Mhb��DM��h�21+� ��������n~�.7P�l��0��S?����j�l��
�'2��Z���ees%Rs��[/��>M�ɱ� �}4�p�#g�ޯ�#�
�S9FZY�?mSӇ?�O�PE� �?-Es��Q�*cb �qV��6�L��m9���6�z=����&,Lhx�ơb�aJ�	8/�v�"���g��� 9�۩��f�w�%31��E�`3�9�wTLt'hU���݈��rb���.j��4����A9"�"���c+�7�k5$�ϑK�F��D�w��4+zi���ٚ�DZA�	�^���Ø�um�y�ʌD�늤�̙�Ǎ������d}#�W[
��ν�ly���9��1f�Ij�X&�����U�C?1|-I��"_�%���wZ�6�s��*����M���5�2p�q��K�T_�c�b���6{�Q�������)e�
/aU��[:3B�a[z�����򟐓#�a�%7��t�����(�Ă\!������JP.�景��g�}��NW�앓�޳���O�Y��@����$9������v�C��ގ����*S��/蛜#9�{���JU�R�i�_�%g�w�'��8�VAy�GG/�86L_?"��V:�����,s������O��M(���WU��@�B0��g��n�Q��eJ��J�B'��r{��A�'A��i��U��:�����Cy�Mn<�-'=M���ت�NqD���m���_*��|�!HҶ�Qe���l�2��Ⱦ/I�b[5�u��T��2hi���C���*:`��yd0�����rC��e��$e�/����8fr�U�.�E[r�m$R*	�RcW#�o'��ʥQ����������ۏMݔ�h>�r+�}uk�"G���d���T�Ѓ2[^��'%���Rה�D�����e7�b��^1dN�[�8m��g��t�SCN#��-����I���2I��Ҟ�'��Θ����v������d�ݓ�]�l��5z]�zfh/^bW�YP��6����ϵ�uuu_���1oG~�P��b�Q~y�v{}�����+jC6�*��F5>��Z�az��J战43j:�S;2�h���i``���2Y���͡s�f�S�h��ȥ��b���vX�H��|��4�ZּՐ��8S���/�Y�i���4�C�I]	��$�ݱEL��}��8���jm�2��d�}���O�ʱ1t�����xu��m,�D�L�@�p�^���8?�C	ų��+"/.+F�r}V���yc�)��UB?��6��>A����+ŋ�VR/��Y�6�W2�����ݡCw7y�>|�|C}�|�O�!����	/V��}�0�O�o/�K͜�-�Q{�7�/��A���9��ٹX����:v_F�<�ǡlw��z�x��]���+��) ���\ZU�t.�|af���\쳨\�Y��y�+��Ǚ�-�n������"���q<Kd����gJV��UWe�C�E� �e]�q����1��:yO�����n���_�q{d����)#�܂fH8�Ȭ�!��6��6Y�B�]�*�q��#j=�!�F��=�ޥ������ ��`7�S�(��CQQ�dׯ�����$�$�Tm�Ú�4=3�6a��lc�}��b`:�\�^ڧQ�ֺd��2S�u�ǝ<���+�Ki����:as�����7�,�+8jq}9�O{���z���l�f�c'��XtL���b�Y3k[���+3? �4�dc7���A�F��o;\xD�v�ӼABzj�G�5RUjnk+��v��UtWަ���v�#$>/�Z�~����OB*�����HY���ڼ���\nJJ
)���G/?����y�U��!�B�a��{�Us���A]�j�vX�;���ni����j��/�C1A"�ԥ��V��U����{������D˪���Դk?v�����7��Aǉ�����3�N�ǆ�VT�B*���2b�Τ������Ǯ}�"�X����`����{����%�0�bwU������w�G;�Pd�ڋ��J����c�(ΰ~t�f���Ž���7����_v������T8�ځ�}�;����.�<�0t���m��*�s����'ϴ�� 2RGE����ia�A�TP�O�?��~�an�T�m�K߱���6��cP��޾�PN���[��]Ʋ�$R#s��[U�{��t��[��n���^;z.����N���j���C�i&%%�l��r���܅Ґ"����wE�������'"�N���-,F�MϞ=��!}ثfmӿha
�8kH�ª�л�xƋ��_g�e��cc���F]���V\Wb�zX-'��5J��ٞ��������{!�ٽ�ϊ�s�pU��^�����=%�Z���+�H�/��H��M�����/,B��s<���l�}dr����|��VwQi�v冽vխ�gF:BO��Q��g��A\�?t�U(7�>A/o#	�վ�ٗ�=8�JY�s��~{޽�q��o�L���%s�G�Z�	^��K����i��r��P�$��i��ǆ؉��W����׌^@��"��1Ӎ�-3%<ۭ쎍RR�ÚY�@�����r1�&��+�J��RE�h`��G�=���U�.�?���W���%y �T�n���O�lWW]��]�'��W7����2��PZ7��\���C	�C�$���c$c��������y�a�������j�6RYY�1騅{���J��z������a�}��/�ɏ�l�N�)�V�t���W���ś[ޛ��D�*zꫯ@���.�/�d{\!��Ϸ�`�󥥘�AUꊽv�Ŋ�M������^��&�%bK��P"�]
�D��,--����J4�����|���\*ب(!�bI��i��܎��f��CR,z8�@���� <�r�.:�����d[Ntۥ1� gd4Y��|lT��ݏ��YN��5Ca�ͳ�� .7W<�x@b�t�U͌E�D����l5�<!�2�̻�˜�h���O+Y�w �жoO��J��r\w����=,{�}>E��[TJ;�C�9ن��~���ݞ�����f&٨��B6(;2���\.��9].x�Tp󷝡V:�)���1%2/.�Rb�A�l�˺=�ȼkęېd��w�xei�(�U��I\I�^��Yv]��5��bG\e��^)7F�����02�.>ƹ�o� �k'�Ge#.,,;��+�ɽ1���%�ȅܺ�;�����ש_���
z�HN.E(��h�p��N[(�fn�xV`s������f2q�6�c�F��x`��H���+�<�I�n�������nBG���;u6e�01!���P�T�Ʌ�K��l���h��=��֍,G�v*;�@�0q����`�Ѣ��!���DtB�m�w�6B��p/�����c���� ��WfyԤ�^��e�{�8Z�T;�_&�q5���?�}��j�����aQ�]�8��� (!"�#���R�)!�4!)(�!� �9��H�(1RC� ���y�������}x73��^k���=3N7��xPMR�7W�=8) �:��Z�8� N`��`��]��w��4���s^?��th��0���{�O9��ӊ"��Ĥ㮘��_�e��q���K��Z%�og������z&L��)1ҍ��FUV��K_��a���LUP���=�ሺL$�[�����z����/�y)G�(^�A�X}��NN?���!oS����4���d����Լw4U�J�����'}�
���Z
ԷM����Z���n���S)+����[LM8i��zq�ߚ�W`�ssM���MՉ�?,��|�9��)�A�b�iŽ�I�U���ƀP�ȼ�1>��!V���H|���$q���5�z�cL�	��c[�����fa��#+c����\駄�����&�Ɍ����!#+�^�	}��8�_vdۉb����!,]5/4T[�Y��N��D�g!5k���������ϣ��̏�ZP!rb�rX�$τ�s*�ӹ7s{>��kM!���Sa�m/�J9!���;�kHaJ(5�� ��`{�{���1�+��7+0����!ꮑMeW>QHH.l9��̘[�-E9Zk/�����b�W���o�-;�T.&[ ^��)i���(�������{�O%�Pm��" �'�r��j��l�6��AOGWP�-ގ���6����n�G�X*Q���D\�]�u��Ed�'�'���;���:�^���F�n���/�M�Z3B�9+�VN�x�V�U@�4�ʹ�AV��SEo՝N�@9*�p~B���39��������n�pF�k\�OM��_rtt:��\0UY�ܽZ�(|�j�V��}����iFQŽ�z+�%h�'��tȪ�=�11.�Hx�Y�����N�4tP��d��5���b���v��w�.�K�yF�����kP��{*�*�α�n�#q�]�����!�����C��XCz�v�\���v��GH�f�4e�ͻ�0�=��r��=�B�qwp�;��d����8�~�r�r�f�?O�h���c��#<����\��no;)**9!�����{�u��Tx[���巠�ǔ�؅Ƚ����{s�V؁��p��4�*��Qjfa�$�M�����T}�`mY�)
��E|#(�������퓗ܕ }K�4���� ���ƹ�r�Y�E.)b�7�꽂�������O'��^�?�T�5��iw�`n���ɠ\]��6�+�
���:��k�V09�����VA�0	����B��=�t��={���}����z��A�A�x3�8�=�����A�ttI�ɉ�#��h�ۿr52���F�ӄ�ZH(XV,�6O4�m��R�{��]=��dUyhSܰ g���ߣ�X��[��N��S���)�{�q�ـ�`�����1[����<5<�=ߣ�����9*+* �-襻�i`��=���R���q{��KTg0)�����£&��kO�<��-K!��?d|-���.����64*����=T�-ju�����ͷgT]c2}4��,�#\l�ԩ���/Eq�+�.�T�*6&?��"B�'<�|��/�a�i�!K��n]���T�߰G�c�O�d�J���L�4��H��\���j!(����D5�"�,[�t�_�j�"3�F��O)�e�o�̯U����v����qZ�ʗ6>��,�Uru�nS�d}�H�����c2�+
5�$�im������Rs��f�9̻�ʿY�Q�Ds�(Vk������b��H��i%�OȲT��[��iB��@U��NŊt���SM�`0��Z��Y����G;�{/SN2��O֬Z�%����D���m��j�DW+y.�������KXn�>=�~��8�{�ׯb]ïBz]7�ߑ�c5�,�{��5�[m4(Mo ��9��b���[�5�>�#(�j��}D3�S���3)�OlZ��~<=dY�ͽ�I�#�.C���C_]��y�"?�O'����`AK�6z�y�|�w
��^�k	�z�PV0�7��r�p?=��5+�nEI�$�g8��=�C�18I�/�M�ס�_~LgaEѿn"���Y�5�X@#Şk���va�����1@�AJ���C�Cc���x�u5���Z�S�qz�V���r>tR�� G�;���
�`��"�N����7 K�e��L�8k���Vٗ��u�KC_X�6{�K�e���X��s���!Tĥr������r����i� 	{�Z��U����Rd�(��QZ���X.z����c'='� އ���R���/|Ò>�����Jג+�|l��ï��)'�9��Z���x�k]�1�E�:@�� �`�J�S�72���@��X����>��gl*u�hg�w��-�}��4�Vt4�'�>������
����uN#������D醾���� �b}Å�b�����2OP�.������ݕۋ�}�{�Q�4u/q�f��Io"י��0P���툝�5U�S�5\EÎn?�x�H����:�0.R&�^Z��He��GT�L���F�E.���T^xV~ڈp���)nzzz��t%eH��[�����O�ڷ��h��W�����[�K����-Yn�(p��� �CK�&%���xQI��P���t@��9:-�D4��!B5t�F�t�l�~�8�EaC=�K�����g�M7PmUz�}|���A�Ɗ���Q/���s�V��y��sQ-���TXg Ƀ�,�!��c>��S�{�ز��b~�W�{�b��>��/���� ����Ɉ�������f�y@��Qn s�����>��_�Rmҏ�j����t�Bq��ɔ@,ͺ�;m4�����x*�$����L�`�RTo���V9�>�m-����9�>��ܝ�0�4J�7�X$$��)'/���~4��ü��p$����AS�oZ���w�e���?tW�}�֯t�	D).2� ]����C����-s�ĵ]�Q��*���N��j��V�̹Oj+�k��h��`p��9���+h�Ҩ���	O.��}��j.=�W�ii�����ޚ�%Уh(&� <cp�5c:�2n�� N�A�"��0Z�G�L���*��O辩H�mlSSI�,�V�x�Z���(
���z��Yo$I��KN���c���sF�k�	���|�&���氵ӕQ��>iz��݅M�FmU����nE,��W�����H�q|�i@�h��4k�8���u�o�U2�h�XYY�	A�`��g��~T�PD���4z
�?�=L�&$bA�GI����]�ܿ��^
Ʈ�AD�Zn.�8��c(���o|B�`4y��un�S�:��t�����T0s�j9>�X��,P#��y0�-?�8H��S7��S���^䞯;p�ݢs|Ş텃n�Z����Հ邏x����LB>�zy�?����V,�%D��V�G�dc<�d�AE��P�t���ISrr��ک�օ��v�������ܣp|t�h���A+��R�/:�N
��uP>2'D�]����,H�N�y�8�������XTX��"��\���j���l�9i�i�L�᫓vMi��d���
 4V��#��3�1��W�!~ݧr��5'���޸���Cxx��ۆ@ۯG���t��t��9�0�7�Bэ��|@�q'''��i�)s񣱸/_@�?�LFb���ht?^}�V)��p�j��_��+��c�N�-�x�)��/�S���^g��P.3�y�5k���R��2��^�%��B{ �4� %Y�=�*��o8Q���r�Թ[��(SN1(>��O�6Z�XZs�`��F�Ζ^շ��X�����	�%"�ܚ�7���� N�k?�5.��~���M�ŷ��<�T�����I���^�P�I��צ��v��nBmg
n��K5��1�X��Y
7���6utZg�M�9��5u����CZ�k�Y�@m��GWO�kuCθ��Ԇm}���2��{F#	@%������l6Z��������̣2��	�a�<�GC���w��vv����Ӷ�!K��)s�9l=T�m��p��p&2����9.����]������d�u ���ʮ���@b���=��+;��B�P1�Z����;�웃r��;����M+����4b}����^��.ÓW @;h�����5<�3���o�}����Z������\�o�ۻ-�4�� �u:r�tr�9Fܖz��	To�}1�V�S�%�_���<����b���
�C�U��c]V��}ҋ� D@�'z��Ժt�sh~�A_Oٗ"x]��2+�I$�X�]�ߓ�5�%*C��-TVh����������w�d�
�{u���Q	�$&X���4Q�JF�^K~ʆr�?>�?�������jBs�]�f� F�ـ�z�(� g/vwdo=k�l�L�S��.&��ATgx �(~�4ou��)�n~�;dI!��8Ȗ�E�(v�ݵ�e_��rl�@ӏy�G���Md~u�mO�]t�wEN-(��;EޞS�Շuǭ���B��� A���H_���JՆ,(�����'����@1
����ǚ���3G�����4�Q�} ��9q�M�X*���e
gsD���3���Ϗ��{�c],�y03�j��s:V�e��6s:��#�1P��R�S��`���BR��,U���uٞ�\ّ�I薟�����*�Uh�
�}���(������S����8�fh|��Xw&�<�w�x���=�}���x:��ϭ>�"��S��y���q�jV����c�}�%s=|J�t�T�C�w%Ùގ���z���:��e����銐k������`���ʆ��fD�+9��ʶ&I���v<�y�,��m�B,�C3�`eo��s���'_���r�>E�Q*� �����?��r��i�:�̊�m:�ￓcu�����M�?��t.'�!t�s �ֻv���Rn�̃���[WM1�$��GU��n�޾ىok5����h�������0`�(�Oυ��`���k�%���!�`ܧ�j�l��F���#�z�gE��6����|��Z_��h���%R[.�	z���)!����"�[&�Д���A\��� C�`_�F�2`�����^G�����O*Myo�������^΅a�>���b�u������;����i��'d��f�}��wh
���癭N��o�Z=wQ���F�2""�f2���EY-U���s}�fs��ո��-Z�����`�����9!5��pYz(J��0��6^g��[��,)�-��d�1WE⾱��N��S�����ӿ�0
fU�j��+�� +�4���z�l{��M��y�>(�Dr��c�=�42=}G�� M��E�>}�he��Ve�JƛjI�]87v�O�������g�����Yx�����#��?W�l={��e�D�)XgT��#�d���FW#��J
)I��􂊘'$D�����H4ltTH�e��^�X�%�����n3�M��w����� 3�j���WP��Sv�_�	\����uBP��1U��U��A��D!��n}?\8 ��^�?����Zw|"I�+�֎�"J�/�i���9If��/��p��b+���(����ː�%��#{u���Y�GX��$qh=����Q'���0' �����Zo�)tܠ�	�ɖ�*�g��w&'dԣ�m��wi)}�&p���1�Uf���2��[���O���9��ͥ"���WS9b6ڻ����z:�v�g������X3�i����p�V�}[6���{�;��������z���1�U�>ch}ܠ�.8��+I��:䴑�d	���%�p↽�yI�\9��.��X�!ws��X;f�;�Y����|0�-i�w*��P|$
2FI�����lA�PH�*��� �7�r^��#U��P�NsrP�ąt9;ɂd��h�����,�Hg>���׫�m�{P��m�a߅������Y�q �xzѷ?�F�EM�>JD�~_`�Sh��c��B���;�׽Q��S��
2N��x��(�2;�.�M�K�L;�_.�#w;t�z����lڇ�1^�mc�{k��&�$�<���#G�n �l���e�|s�>��ۨt�w?=9ޜ�Tb��l{}�6�_	��U�k�h_�B�CJL���Q0�i5_�d�wH"�J�Y�k�&W7:��:��g�og��YШ�ڮ(??�nt2�����{��T�$�dP��֚������Td1�{ �L�0�GE�\f[�g��Rn,VH��:�!LΈ�D�]_ULL,nb�����j	]���Md�Dg����;4�O�q �{�)¦��;;;��]yY�B��6�qU�G�3�2)6�ç�}	�FcS)Y_^Rc��뗽�%GR��6i�մ�Pye�"�3�.�E����P+V"����^K���������ɱ�
 �ex����;�vO��.�Gzt�l-��)�����X|�"�-V�V���|V̩���������R���%�j�����)�'�񂕭��@��=a��Z��+�&����?������	H6��,[�[��d]���h�OLL�ߺu��y���9�_�#߅������*�<v-7��^��jC�3��(n�e�k�w6�N5����͒:��8�XN�φƈ~�wj_7��LȮ�Έ�]�>ݲ�v��K�w<��`�(MP������\TG�2U��5f����QTB���%��B��H�m�t$^p�������_�06���R�Y�����gf����J/<�qS��Q��rM	��/F���4�B_���+���xu��p�]@I��՗��ȯ�o@�RA7a�C?��#p�.����kc���>��>Z)�Ge+�2|ɡ������:tC�')ULg�T�@{G`����{Q�<@ ���6�T�� ��R��v{��oB�-�3>S���s$�,Um��4�:��+b�C�B�nwu�/Ե
C�% ���j��|��g�G���L�}V�
�e�l&;; �-���
ލZ�������D����zIƝ�|�d� �||�#Ŵ3��qY���������-Z�M9�� eF+-v��[��Q�G��(�Ł��z�����|���M�>��|or��W�f�،xW����զ���D��0�S�A����lS o��}�V��mٛ��b0��8Dk��C JH�<A#AQ�S��U� ����8��>u!n�ۢ���7�4����|W�i�t�\;&�w[�!���*v�wp�x��޼{��Y�/�g�:N�s
��=��$&���f���IK�������ӳFG)�Q*�c�%�ˇ. BM�?m�����*�GG$�Tw��o��q�0����M��ˢe�ư����3��������ΖTj��6+3R5�RϔfP���74ƶ���0j�W�f):���R��S���vJY��3�@��nQqޘ �ݛ��tYv�77�y�����[|�e�IZ��U� _X�e\i\���$�\gyi��I�r\��ӿk'�%vyj���S����C�W��֑��R9�a��|��K�΋�Y�RV������c\]�n�@�I1���D�e${l>+�'�d�4�_����B�-�;飤t�D��ؓA+���o"�̠��V��ר�m���nj�]�nl�k,�P �7z	��H��Ho\=B����h��Gbw��l!���V�~�s2��6���ۻ��D�Yo�p0y���+[l�T�
|N1��'ίѦЋ*;��xD�u�-�'Ľ��Yht�]U�t ��@��������o�8z�!�IF��:i<$�Sq�4�9��ʱd��a[�
�x�#<_�%�F=�zp��̭��:��@�^��%�~
�m�[�ō����N���Q�L2r�MD��yN�Vd���|@�,��?�ip�W��%�o3>��C��L�*~�D�Tc��9��!��+vd%<��O��;.b�$�D���3�<q�����Sf͍^�������W���k��"D�~��VoKO=��z���B��#�='�H`�q/
�Q��Q���Q�A�`��v3?j}���h���Y,�b�KW��������gP�$YL7�������ۣ��,
�i���w�C��\^���,��qf(�T�xP����]{F]����*��1��XQT�?i��ʭƲA B�-n
;d.O>�*�	�@�Տgp�+Y�銁\K\m6>�Q���g���ۧw�^���4̄]{3����:@+1���r��i��>Bt�����f�I@ʌt�Y��a:�Z$˳��c�]D<��g���i
�6����Z��W�F1C�R�6*ߖN�3�.�P-�?!W�z�`�Ü�ʽ�Fu^`$����&�ʃti_��6����`ؕ�Z9�7+ *3��X�����HU<����X� ZQ	U�ӳl<.�{��$-��������ob�L��S<���VΒ^�YTg�N��;�ZO�c�ם%�>�i�*aľP�)��5�4�&n�<�W'�!p��A�)8�gmm]b�8/4(��o����b:�td�W	[~�Y$��������9(�TJ~��I�iPYub�u�6Ӡ�(Í�Wt�@r3�6:�kw��.A���'0���sB���9��m	�Xn�t����R��Ԉ�(�uzsf�,o�:�u��Z\�\���Zْ����!��V�z��©�.d���S,0f}ԥ7���^����~���i��5�p�#c�Z����(#U�AF��t���K�`�h
���8�]�c�k�߄�):�4����q�F�`����i27#�����Ɋ�PضG��P.DbtHH���2>�UK1½LĎka�~�t�UV�]��3O�q�sy8E�߽=�+`9�����!��͟L�Y�ڧ������q!VrZ���M1r��oM���i`�+J�]%�5���}�� �ԃpf``�FH␄6p�]-���23���Hw�~5�������v�V��$�x��A|�L�-�l�Ь�wn:�b�w�e.(X����}b��}���X|�wW,7���w��[�}�{���5�*�g\(g�E��>!B/��o����/���Xڮ��]�DPzw_8@��>Kx�&�Ѧ"K6���/��@�K���ó��X��)��獣:�#,�1,��j����;��)(���MJ�����uP�7�[T4@��Ï���^~ڦ�S��Å�����b��(Mb���~8z��s[�ʬ�{���S�4xzt�ƫ�=թw���Q�w�����콷;a��5a]q�`�]�VlOG�2���%145���{4u���S�b�Q�Du�jar\o�H�8��C58t����"ˬH$o%�{4sB�b�J�*��cH�u|�y�F�Vc��e/� ���V+fb��ݕ aW;[Gu��h�z��G���y	��	��&i�ӊ fr ���ߌ8[x����[X�	NîsN`��W"Ia-�tQﯶ=�\�M1ٺ�[ӳ����ݬ���T�A>��*�mur"����oPL�U!�cn	�s��~ybC�����Bǎ5/�o����v-�����L=c����e�`eȇ��[�z�l��ě����u�fn�~٧a�%�f�J~c�_�q��0���>��SVt���P�2�Tq�Lq�P��?��^�#K��=ZsI*�v
R/k�~���qB�;N��������1r��.�͚��)^&@���P�x:�p9�@��R���}ԫ�D�ymIF�BL��������RǕ�d� �J�5֥��̹{����I��{�v%�\��eo�j��r���a*�`�\V�
t!_6����j���ԯ������O���l��X�Gh�R�1���R'��
6��[�n�p��<#F�N6W�xe��7����C��NĄ�I[���X�XB�몰�5ٞh4����R�=��V�����$�ɗ*�����K']�=��=���My�*���/ONV9f1I�����c�o�K�*�>}���/�|0��X�K��
6������5��#U���rs+�8�E��B,��֏��J�9���"(ب�۫֫�L/&�w~f	���|��U��kK';E
#��t����e@�skDv��'�F�}����o��/&�B>��5�A��1�oҳ��p�/��{�����?��+<�'A[5:����D�<���]b;㥽��	yV������{E���JQ�e	y��w8|}oW�2@�c
��[��x8�k�N\*���!Ʊ�7iY�����_ã/���?��qh�栩}��n�����.�{�I"t����?���ɉ����4�?�B�b:��������c�y�R%����2�M�oS����/�\�p9�p�I�b�}]�I�3�!���8�nG���Q���޻k���LU%˾��߭6*����}+4�'�zX	ò�b�[���k�QTa���8��i�#����7Eu,o��� +mP���]���,��Y�m����c��w�:�����#~r#<j,!�j�t�������*��8���Y6Ҽ��$OeP�@��<<r�M����c�AwM{�/G���#3U�ķKy��<^�p���Ehd<�3"�죴�u�E*V�������� ���}b�;���M��Q2�s�ɋrpD��h]�s�8��wb&f��_u�JM�W���3��5�P4�tQ���J��=���kϱ�٭g�nE.�-ּ�P_mʻ�I�"�M�e��Bn��(��w�	��Υ��c�����$�7*��F>�\����Ɖ	�)�x9�͌&m�R3�] �����H��,Y�r���w{8������zo��3\;�)2go���:.�j��D`��2�{a�w�r��Lets�r���rw���V@�z��y�y#�C��5�bػ\����x�����2���2M�E	���ҙ�hYݱ���eާ^c�LBJW�f��t�׷��M�m3���|4/�qg꜏���v0��n����*Z�1^�B�E��Ñ�MW��(��ʿ?�Vv����F�F�(V�V�`_U*�����;��1J��^*��+y���=��kq�-ԯ1툸L~�W¹8V���)��0$`3Y�Vl�>m��ag#r!X����~i�g�Wٽ�����/��HI��9����7��Ŷ)�~U�O�61RL�}X��u�I%��2kٴ��R���\:��b��_�Ӯ˓��T�9��O"S��'����Zy����?ڿ�˭���u�*'�9)$�%Y��J
��f�D�������K��"�H�e=@���z��×�$ױ���E�_�3]\�n�ccl[=jQr���Y�ȰM�]��R�,�.��ׄ������G
![�%+N^��/D_��A�&W`P��W�&<3/��L�<~协�F�K� s� d˾*��Lu����<�~����K�Ry=��~+������ྀ���Ƀ�k�8�W��>>R@�O��rY	[�/t�3��#�!�9=Rnyh�X�� :^��bf'Y�M`%�mkWq&�ѹ�===Ɨ�Ih�ã��G��������c��o(wAo�l���3';U�������Nʓ`�(r�i�4'��K
w�,�IA���(4h{�� �!��>*�z"j�.��.�0Y�覇[eƍ�.�ׯ_�v�E�.�m1+���p0���,�Xn�e����98Ȼ�Y�	����vHe@&��6���]|��v��y(�����DPB)�"?�a�h���,���?�:�A!�7�s��5�%�?W���K��W�O�0�V�x{�s�gϞ��A���4��}��]=����K2�nCVV�RY����H, �����h)��.�i��L�G�k�[���?@@�ܓ;l�z�R�����2r'/.Y�[O�����aQJ^��x��z>E�
y��z�">�:�q�5}Û��4[�\۫r�[�?�<ݲX��s7���H;7�gg�S��k�O���g��4y��W$�i?~�~�G�ҫ��$��u�D��[�%��<�<�<�I����Tv���!�������#@~�DE����Гp�s坹���<�V	{�:h&���:� �̜ѓy0_�s�lO���Ԯ7����	^��A�6���$��[�+�9P�!��k�5ZN�%�y�I��{Ue���2�� zE�ܕ�������	ѽ"��%���9���O{y,���k~TT��t|S���ɕ�Ҭ�����	R*8���Z�����	�3������^̉H��s;,ē-i���V�{��@�b\��Uz��وu���.�t)3�T�-@B(��\������4���M>'� F�/_���Z�@��J���-�LU���j�I�y�� 'i��0�Y!Ǚ�����v���[��!������|?e|�@U�B���7���ڂ:���VS�UY�~+��)�1�o����d1]���9ܳ窇�F?�q��2]�["~��犔x
Y�N?�� �����}B-�Ғ0�����'zc?��H?[9]br���,�"�P>�7{��_J�C �aH%�k^�}�׌��T~�۟�Id�f���)I�3�//x3��gExX9��^��s��ś�
T�U�/Ɨ ��~ދ����M�c��w�mg���5���c��x�	��l�%M�s�#��w츂��rK�{��n�H9����|�GRL50��;ܖ��Ol��]��Cڼ}�ɷ�p�������gv^dv5ΫU ������7E�r�G�������]�\���E��0-��PE�k�o3n�p>�$m���|�P�#�m_ͤ�m�< o7���O��(7��W��u;1��'G�Ie��Z��更`��)��|����%��W�e2�O6q��A^�p�.�6(�W��ܙ��|����[��Õ������Oo5Z��?�K-v�ظ�2�t�a�Bܗh�t�]���}�"�/y�vg���� �v�/*����k��3��zSh�L��*t����y��]O���Ϭ��q-��$��2�(��:�T��ɋ�`�we��"���0D��9ي�1]}	}bG�n��A*B�L��>�ΰ���,�׎��$5B�+���U均�1�>׎^�:�AO��L~P�L�C����/A_V��ƪ�W��0*���U2����fed@�~������はM�3���2`$�`�������Ŧ#t5�fc�~�W���ϧ������L��)V�<�%BS&v!�����Z�z��yf��������=%ѝ�t)��!��b��;���X9�,���z����R0R�5�U�k�'���|'�	��C���a����h����w�n^��eM��<9>���}�����M���aA ���H��|�s�3u���s.Nh���u�)x��D��yO�]&� ��

*|��	�AŮ��\<�؋>B_��ZLL�V/�,����*������|����1�5Q�#��IF���S����P=��o� Eb��+�+�|�,���n����ԍdD����c�ԁ���;�]����y*c9*S�X�]�*S�%��d(�2ce��R^NfU4QYZZb6[�Ӏ����U:n����go�.�=��6x��r@�=_��g��CO_�*�Q�g`����B�X۟H�[ڜ	kfd�@ީrǂ�w��r��8$[��K.`	c����Du���_HE�^<�i�fӉ�\Q�0��Dc[��Z�`����:L���W\���Z���Iz�CɼqϏC+��M�>ۂ����؁�Ne�j"Ǻf�#񚆞�Å���nk)ޢ���Px����hd���Y��~�'��r�^����<��l�V�5�U.EPB Mm��%�o�~C��A:#B�
�P�������0�_��ua�@� �d���
���QRd���%�3��'n�s�8]K�T�0���W�OX6�I���6ѹ=������hټh�I��KS�9|�<#�3hN�:Z嘃��|� ذ(R꼪�]���o����bF ꖗ[��.��+x�Ho��|�U-�V�+��.�d ���F��� �	�#A[SR�g����@U�!���\�H1Iv�ho-��!�i@@L�k�U�<��8�J��n/��[�c�ECx���  �����WJ��������X�cz��O8�#��-6U�@V��뫶����|P���y#��t�>�����X�3ˬ�uy\5�\��J)QH��lwo��,�P~,��χ�|���&��(qIO����uN����m�Ήr�v�r�>}Ϯ���!0D�9��DhFƛ�������0�!�V�����/�{{��.�{M`aaFc[���MVe� �4�=�V'l�]\{����w ���E��t�楿/:j�d0���*��Ց�8?]�� �c]�&��ҺB�n1L����y�[ރ�]�Lx���tжŰ�-��pee%�`�!�I0�����,��k��1@���;ڿqM�K�����C���8�4I?��L���� �� �_�w��n� ��9n*�oN:*׼���k�)�չo��>���1I���d��������ggk"@^�	̯�7S5]1��.�k�]�������gN�O���gĄ;���^���
 G�bkGE�f�
�?D�"�&@ُ:ۉ��më,t�c̀&������� q��T%����X�ݭK��n���LT�O��jyFCL:�|�]7��|UC�q���St�b ��ul��j���z������y6�:
�x����E�?��2k���
'l}� �Y�26Ӊ�|���?���Sv�t<T1�HU5h�-�ߋ�a<��[��T[������y7��S���y�H����4)׸����8��j��,�gI�%N�2��1F6����9��Kt��t�.��Ժ:�(Ŏ
� 9��[!_�7Lw!W�T�$���^|����߃���Ͷ;3��J�u�$ 5����Ą�>��ޔ����@���� =�ǭ���RU� ��QT�|���	�T<T�JO��m/C-��d���f�'���z���Y�ߢ�C-��d	�G���#��˔�hDDL[�Ug����,��~Wױ����?]�2#K���2��Ʃ]Ȫ�f�ɝ��)��&�M����,U�e�#���]5G>RH�V��P����|����*l��=��U��� )/�W�q��]�0�oh9���� R8���^���b���y�)���/h��r\Q�f�pG�'�,2ml��=*Ma���m������
A��d,,�r;���#��~6������(�˰�)��]&������d�|�G�ʽ�Y ���{3Egz3-l˯H�v��+�K-�w���b���(-�u�A!*�D���m�{`�1�u���1wP���W���r��'~V�P3�F����<7�O���,���T�H챫܏f��{&�E58������Cp�ſ�-(�D��w�G��S<�E�j�5����I	ob(B�����RV삢e�o���B`RB�`�^]%V�H	 _>�m�����͛�v�kv��u���h��j8��\�YH���Y���-�������CU�>�TVT��j����l�w��*?H��>��L=����+�"p�����>����p���Ϟb�^ �%�>{���0�۫��\���۴�%�2�#@�0��C%�j�������J�M^p�me'�����/����'��F��bzI$�6xZ��������	p�����q�M�+Z=l�ʄ�c�<X���.�$U��r��+�����@�L�����
@�F��Dr�^RwS�[])8rw�NT+{4hQ웛]<���n� ��z�}�2�ϳ!�l� ��$���K
	�9p�%���8\��(g�7b*{�e?���tL���u�*䴆�d%p9�����;���\�o{�vhӔhH�
�˴�ֳ3�(�F.9�z��M.Sf��s~O��Z��?�it��J=[�6�]�~-|�f��v�>��o��%nb:J�{{���/��\���%n�Z����w���?T��9�;#��z�9�ve>R�y@l���g�˿��<ff���t;�{RL'Q��$��E$t��?#������ȹ�rP��RƂ���SȊ�>�+��+R;5J A#4��1㔏�5w�~+�]�=Z�em�8$��z1��X4]���b�8Q��d#(B�t���3�S�����v����s��4<vì�BЏ�N�.�jҟ����6��Q��ܯ�4Ⱥtt��;�.�\�ڭЕ����J��=xHb� �����c� ��J��@����b�w�ݨ�u��7<�+��dM}Q-c�~8�	�r�aTT�z����Ԛ�����̃�)	��~��l�L	-���S��� �ާ�w�S���������M�<X ��Ja1RIE��-�k(�5XZز�|�O�K�����dR��] )� R�ja�f�)��Eqٛ�N��c]qm�n~)�P���(}�ݸ�D����÷�+�z>�P���_X�KS=�M�6�fN�A1�j�l�@+�)�4X�kkk��v̒D�L��������3��:u@���nzk��צ�B�x4 �ǘu| c�)�T< �%%tC�8󉎰#����4��5�)�G�s���9��&b$C�BF=vC� ���2�_���U#��[�Y�JG��@e�������yOpƣ{o}a��a�u��"�:��L@ ����U�ޑS9��Gυ$���4�����3�,��X��1����~�Zu:@�6��#�

z6v����a�$;V����AL�ݲ��-{���B�˿9���)�u�K��A%`�eBi�p�H��� 곲�z�c��
"1ו M\�����<*J�\i���$��AǨ�x������dПw���V@�͡��!`:8>Ξ�Q𛮙v�¢�񵍍F��'�:�?�#@�蝴���đĉΑϹ��Rl�=ޫ�)�${�<��<�����b��? ��If|V5��?V54,b���
�����l��e�ʌ[u�K���I7y�s�Z�b����i��7-��PB���C|�lD^���|̍����OFhD�h1�@�H*�%U��/.�Ł�4b
���������V�@ʬz|�	���N��{C�@��Z��'4P�7��pH�
R�� �>=�-�d�n�Z}?v�/��,dYo�f�2��&�)�y)/2���0:�2�ӿ~�2���}C_V/��?�.��R��K�����Y�3��{aw���9�j,_ߣ��Bw<��\>��W��E �`�,Xﻓ�v���.�N�[�1�����������X���)t�sX�0h=�#�L���������OD?�hFn) �Zʭ���&5u?/{3/�p�	083�aT�#&vqPR� )q_?��m�`�iH�<����*ya�jߺ��8`)���H�=ʀ�7��� ���&A;��,4[? q�R�;�7���o~S�.U��`��Q������o��
�K��t
�
�\i�ːJ �qe)a=���5�����&�K��j g�2S���/~(wk�p��@�v��
��%�!����a�n^ �T@�%Sd�^�f���s^	C%�?Wa<�|�j�ov�Aӑ��8c\�Z�9v�-�X�̺�PƆ�R�0%��8U��{w��П�F�b����0�����p#IhE����/JHI��b�+l��� ��
�t��T����8��[P��LU/b�KR�C1i�X�&��}Ƌ��)��w�a�a돤6�F��Ԥ#���xu�x�v�k�r3y�{������$+�X�1�c�jڇ5=�6�r��t}	4�mԶ���@B�B�P�y.S"�p����<dh"N$3!�1T8f*���9�c���?�8�����[�]�w����}�{_�������K�2CU�����b�d���-L�0�^]��Ax��庩S�'�!J ��J	$�Z'��'b�5p��k:@�ɣ��B�+~]�Y�4�J�x��c �!�u�T/���c�������A������C&3�n0������rO���x�t~��G�%[�.,�#j�]8�t|��٤r�?��ʉc�>��:ـ��w,��<A@X#���>��_�r`���w�	���Ue�F�څP�i��W�U��?��'��N%�D\!A���|��5)2���`���*wSA>���~�4�	bS��N���C�A����T�+_N,mSgh'��q��FM䩼���a\~W�a�_��ۉ�������J����"��;�9g�vaq<O�4uͩl��bl�mhb"tCF��{�Lj�c-,,h��3XsTw���"C���_��r�Rg�����Գ��?��V�Fi@z{��}y��,��f��ͩ�r5ޘ'ŦXRA���%�sl۵K u�vV���I�"�¥q���O��V�噀d��:ϔ�/C8U�f�ѧܪ7�Sf=�11������j3�N���k��8��C�6
i�R��BA�r�^�:O��RQ�!���q�i ���B�k��!��@8x�a?m@ �	���K*@AH%�U͖"\�FV�ѨI�̄��B�`��w���D����W�	�=g|J��U�;����{�_C)���W�`7D�|��Kp��{tQ�!�9$34�5{�mG���5�os�RO��.�#��Z�3��D������	t�aӧyy$ʄ
p/����b^l��L
{�/t�P���S�}4�����מ8�ckX���)�Z�Br~>�S�K�kC��4ueF��j��+-�8�O��;ߺ��@:�z���ݻ����V[N�i�I��#]����LϨ�CsQ���f�*��;���f~��N逺&�V^H��D�Kp`�>d_���_�7�Ib�b���-x
� �h+�E�9H�.�iE݁@ɻ��Gǻ	q�E���(Βêt�/,��O��G��Mg\�>��}'O=��UR���3f�S|322���Z�S+^0��(��ڴ�oP��$:�M�ģ�	V*e �)�@��,��`��|djsF&~�#��\b)6z�ށ����꾩�v�A�4�<mp@�o��(5�vAE=� ���r��Ⱦ��3㝂(;����w��hI ��u�C��rL��,v��� o�
�=A8�>�j����M���	R��ڬ�f�*^�+V)C���)X�rH�q�	�����| J5�Ρ�W�*fg��P��R����Q^����Ry��qq���r�!��lV���O+;�d�$�"��5�Z�o��~$�hTѓ�Mf.\dW}�@p$f��Zd�W�g3߸޺pjh��b2tZ���;d��+���� GpvnAv�'�iC:�z�<vL�Y���;��iL�3����wA�ֺ�/Vw��2�W-�Jҹ.I�����`n�}�Էu<�	��2�S��3�/��S�jQ�����ʭ���_�(�50�27#H���4�ԉCj]*xd��=�N�qZ^S�(� �6�� ���%#i�q�JS\A#�Nr�BpW)�4�K�֥W�/4����4Vݤ�޶��?�Cc�W�;�\b���ٯ9��ߡ�ڋ�%-�����/�P@�3��6���™ѵ�i7v�IާCv1|se��r��x�q�ImE[������;�1Aq��I"j�u,Q���U�@�T��3?qi�5��Zj���y��ẓ�-���٨ �U������v�������ƥ7k�2f�ب��MG�S�~�E��'�}O�Hu��pJ��%g� } 2��w�1`�X���������¯yrW�+#%^䨦p![��CۈWc:c�빶�ըٴ�	t~_�шw��A���u*Rh����>�)�Z��[���E9)Γ�>={�������G�O�n/\_1�^�Y�!��KA���������N��gk����iyb��o�(�?@m"���O1ہ������Z�lǆ�7�}X�GCL��<��Ŝ*�*�DKvp�m���zy�X�xj���z�"��z��66619iF8zK{�a���V���G�P��=�2�ۻ3D�	t�`�A�;��S:k���~<�6+��sD Q�WB!���])ר�J�$�ɒ8n�zh���a(2���P�:�����;���(�Ly������R��G�5�G˖U���)[(k�`�c�.���?���ϯ��퇲/�\�hK��/���6�?��2Z�U ��������g���O�5)�����C�^u�V�x5���I91t�>y�$G�g�M�o�}# ��P��n�!�S���as�O-i���l��S�C
4#����J-��o���!���>�s�[	���"�s�o4��K=sV��6v�?{z|���]��w�;'����xļƬ���[��83	��)�s�����N'XS��*ʊi����n=�cO�d��-{�#3��6R�6��.}�YB�^�w��&b���0�Y�B��Zf��<���:7$G�|��+�k���Q�eYԭ]���t��?ud<
˒��XM�	W�{�8�����讆ٿg�0n��5�q0�N��z��X�w�=�r5�7I?�+�������G�6�1f�;(��A	���AY�@"���_�7iJ�|PypY�Ro_���G��2�8}Ӯ����`��8����H�vܔ�
��k+M3����� �m��L�E`L��A����7��P��9����/u���-��]���{)���p�SF~ڬ�aR�Aμ"�^�T/�^��q�qt?��ha�9Gݣya�v���q�р�C���鳡꛳��,g:%�^�Rלh�����1�4	����|�(e�p��7v���i!��S�y����5�}��;�l��[����>Fh�Yխ���u���fN�	�U0'����>{+-&-���T޼X�n�蔴��I��<
�����8�O��/�HD8��Q�Zk��2c��/��������0?��%� ��wM�fB|��*մK�g@���{�	�:�RJ;1��?)	��u����<Y��#k���s��;�@��!Gai������9`�V�������L��ʣ�#`����[P��O֙9-�Ͽګ\"��T�����N u����U��֝W�.���N�L�J��1R��y"\ �9���*�W���9���cf߮*�Z����,pڞjF��������τ���2��k�!��i�����߸ ��W&��c|�@�U͟RQ~��T��1��l�Yq�+Ρ����҅�Ҟ{6}���x�������t���|E؄�+w�L��DQ^�?Z?F�)zX��m�5揰hp�6��:��|e�*�b�j��[cmQ��R�I)����y���Bâ���~�"#no�=^�
4c?"���;���3��C����7��0u
v�}�Dg���@�r��p��vw̤%��6c|t�Y�R��2J�Ϗ���S=99�ő9�"���}��吹˥?�\� �9/V���KH@h����\��5j�܏М@Z�@?G�R��+���Ԣ?o4�ff)e`�Cv o�F.�h�*�T�����J��t|���@BL�~�/P�f�����hVZ��ly�V�_�;O(��̋j7�dk��`���N0J���;~'n��ḨG���3����)��O+���=ڪ��ѧ��G��Xo+/b�	�.�m�OD��Rr�;E��؆O`o>q�Έ`�Nr����%�����qo�E���j��Ɛ>m�B���C��3.,J\ s�7���x�N���E��w�V���T$Jt�p�ڀ/��{*�������^F��<�+hx�$�9��E3���a�d<�ʆ����e�B[o��D�Ѯ�����ֲ���ן6/jTF���2��Og��~xU�_58��e݂�ލ����F��ٖ��y�7,^#�����Nk��(֞"����026���[]���D0~�(�<�S���A�z���@�{(�uP]���@)���JN}�L[�!̚

O�.?�S2p2�$KǄ7*	���K��$��,)�Y�W�;R
@f>5�n{��}��+מ�
�#��T�椸lǉ�����1w^{ 3;4�
t�9����$z��?��Uԭ��՚�����L[�v�_�VV|6T�G�&�8�K���{�CԓE���c+ ���\}�������Q�8���*z���T�W���:_]����~&$C�o�v�Ģ��d�4fd�T���o�dpl�3�K�Ɉ�~����N�_  o)�������K�	�g��KJEQ���<˫ �����M�=�+���hk)<�'���g�׶�$�gk��,S�s[��!������w3[�&TI�h�*��&�y<=#$eY�F?�L]�/�':q
��b���ۿ�!ǊXo�s��k7]�0(�?�q;3�Ϊ9��.��=f\Ą���V��,d�jm
 ���1f�I�����;52=Fwg� C�/�Cc3���C�H�UB�#@л�ol����֌k�\�9�Ty/����ܭ�,��B
͑�z(|Y�R��\uBc��GE
�<F�(�&��*�eۯф�j9e$��$�sGz�K�/����	Ks����՚_�Nb��	bN��%'���Ӣ.O�߹��!��kʖ�=��I������~	6Z1���ABq�Y7��������5"DBO�ӳ"�����S�ІOKa�31c�c��$ �Hٗ>BX�?�v��+�?��Z��EF5�"E �z�m3>��Ψo1�?�u!��m�[�lqv�l�]�ym��"�4�`�E&���X=�0w��� �X1����
YGaS7������?[�r@N��Tf��(�oI�ǫ̫�o�f32�2�_�xj�����6ѓ#����⫴0+
>!���"D�T������f:A�G��ޖX����ݧG���\�����S�)�b��9̙���o[�E���Ƙ%3 7��1d�)))1L�66��Pby���h�Q�ؘ���c�tAT����C��&�:>WT+[t�˫�G�^�@����.?��0;��������?ߚ����P� �1K�9@�Ҝ���o-�&�p&H;R�&N���UuҨ��1�]�� &UrPt���Y[ �w��4�����2���2�/(�������+���c�������F���^��a�r�C,��
����13s�T��TZ[�����#��M�D���Q�����vv������g�^��?K���du3�����#�[4Dr���%w��,bG�����I�~�=�ؗ�G
H�9��C��|���r+4J-{y��.�B7L�����6u�Zz�ˈk���l|o~<~-��t�����?�3L�5���D�n�uZ������N��k��u;�z��V`߳��R:g��4 ��1!��j����{�N��6�$U�����Cv�m �������� ]�/�Bad)��V���d�w���*r��*�M���1�v�m���% ���Uk����`��&T�%z��M��G�I�fF��&�x^X8�y���Zr��x\>hr�*�$�{TW�R5��3�f��f!"E��$�Ǳ�#c��(�2�SBC�$<�������`�%�L~yjw�$:7J���5Vi4a������m�uVG�O�z�̨�'�Rs@̂D�.<�H�XSzy�����f���2o�a�Σ�+���J�6ݖY*�%_�D�D�4�2���O��%�e�lq/����r�����S�k�M7{?�`+��.���n�3�w��oaDX��Ǵr�V���ܦH%y�x5x�P;���`��766Z-��Wl��s�?�Mϸ ��D��q����C�>j���/60���in,z�߽��3U�d�2�<}�f&C�)�����5=VBfH��k>F> 80�j��	}���@T�#�u��J�Y�3!�@�!,�Յ��c�>'�{�Mh|eQUzW�$o�5)QM0A��O����� �=�m�_��v����u��p� Z0�����h�~���6:��_�(Q8��n�Ɔ ��)��Dɺ�]9��ok���FS��mӓ~�Wrd�c�Z�0�g��s���g�v�e#r�Y�a�v�ٍ��L$ҐE)���}H2�];����\���޿d��hn�E�Ѩ�UW���Fj`��c��$Lz��ww�*b����2�Wͱ3$9�.���+���Ϯ�[�QK�iyzbZ�/�:.
_S�^��h9��P>��X�3�}r�<��8}��G\	&��1K$K���s�y�?���'�l���9gAV�:)�-m���کKScR>g��#��)�,�<߭O���pJwB~Iq�rAQy�t{���;
=���<�㼯Z₸��D�ZFUzdǭ˃�Y�<����j�w�WȲγd!\�g%��v��SMd|��Γ׬G���x���,�%������Qg��IO��N!:��H�-�peͰ��	#$�R�K����b����[A���j
��_.���Į��+Czb�R1`|^ '��,yh�h]((,{A!��49X@��C|������y|�;u�oE�~-��8fǱ�OT���^���������"�q\^��x/����{�lc�Vg&���5�p����5b��y��Z�W��Jg[���3kUSo�L�pHK�'{���O��T5�G����!��N�E�9^�q�R��TM��kB����C�W�	cX���g����r�Z���
�p�۳�s�y��(������$n��gJ��>]�G�B&|�QVNY�P�,��R�ڛiF·�痆��s:��]Nvx�T�ѫ6Ad���ס}����ף�s���}�fr>w�/��u��� �5R�l�3�-D�L����'WkiT�+;bBG�=�3����p��=/�#��D(4�9�5�_�;sV��o�����O�a!wO9���޽��[+�f���M�`���[p�X=�Te����Gll�afdD��"�ѱ�7N��E_S�q"�������v@r�oU�V��Y�o˧C���B$^?W�"��^��.�m�=9���j�.�W5őJ$���:΍�no�]������lF�OFi?���a-�-3�$ ��Gaj2��CB|mI3TH���_ɇ�^"��H��{�n���G�����O��A���m�Q�����P��M�odYHp��g�\�Z��D!��,�2�I����H!���?Q�Q�*-�m�w`�1��5�Ͽ{�տ����E�x�v��I���H�(4�NfS��9+d�nIi<K�.���f>�ʏ��G�1�#��A��Q���O�����8j�y诵}!'}��)�g���X#D��H$wN�����T�!�kܤ��&G5�er��&+�� ��>Z#� `r8�S;�.W���o���Ӝ)&k2� ���z�&XCT�_�B�J�H]�m7k���Exݼ�"�������\3�V�Q.��Xٲ}���I:w��Ї.3_U����$�|�w!���
pʿ���O�[}5ꅢ27k|�z�ȗA�ƪ��q��b�|�L9Iq.碆�}rr��4����}��$l���Qy�(*K,%к*�a�ڨv� �E�s��H��PW�SP4%k�5�Du�<��Yw�xqRcc/H냙��F�7]�񪫫�Ix:/���kh�S���8>Q|���>�z���+�d⽾�V�ȟFvy+Yon��@���g2_�j��M��g9��[�[.}�u���'"&�O�V����n2x��1r��e����u7!r<��3�����d��~/7���hV}�`�$�����!�Nr��*��#�����iU'
|X�M".�B%���ǆ?�29�+;J�[�aN� �G����dY�D<S����{�yr�L��'� �ld�T�Ϙ�o���T|�ݣ*þ����9K���@GI���3*H�5�Xf1�F�x�mb�v|�B�@@5�>�Z�D]�����r�3���q24�&��\{$p���[�$��IU�#��̷��m��(q�A�r�L��ީ��Nb0e�R���Jm�RH	+98a#{Vj��v s �ǈ��\lHTNn�|]=�2y{��0��쒁�E{5|щG��������*8��b�bڞ"W|f?�P�/"E�mX�Y�S�L���T��J�J�$�-���6�l�;��q�� h*�B���9C����z�U�fԸ2s
/�[
�C��Z�'ʤ9�{�u�s|��f\�ڴ�µ��	5U����V*�	���]c2 ��EB�Y��@{����X/�Y}�9�.؃��1|�8Y��f�f���h��ѷ:�4R�����9զ�h��B�؈0��K��L�s]Fو<���$��v���S,����X���uaa��Ԓ�v��1�F�[A
�L��N��2[�a���͗f:_n�([�1��p 9K|���܊
�p��<����:���݃D#�dL��#.�@�w�������4�zY'�@Q3��- !��\|�A��Y��_����Q�4᫷�	c~3gǍ��M���h��@�ن�� ?����fF�c?����邡k|
�ʄ���S�y�ACuu��K��3�E��P����e���������$�2I�\T�_9φ7���I�2u�TV0��V&�rLi��&��Bz)L�b?l���'k��'dyܱ��)�9hیJN�&�>o��
|��m�a����B�\k���i��j:�>�ʀ(���^�R�bS���,���a�|hh"p@����?����sO�e(�A:E��:?�V�\�!)�-�pE�l�!����r��h�
�4s��m<􌿖k�5������,�<�9XT�X#0�b�����f�&����rvalk��
:�O�:�q�4�3�! ߌc�믵����|Gǿ W5��!�%���S��XJB����q
JA��q���j���B Jo�O���V�5��a���1����K�Pb������Fµm�&����\N>_PoU�������G��C|{��"�^�D��۳����P��P�xU.��F_�#O>�.���q����"cO�������� �u����}�RŜ,Bʖ׷_�D��O�y~!��S{��T'�w�mŶ���LT=Q���Z�z�:�sts����4��5 F�W��aj|�Ȟ��'�O��F$��E�sf8Y:��`n妷,��nL!8����g�?'��¹�z��,u�u���g�n�n����7T��Ӆ��x���<�xU~6t��^��g�^)���Mr�CIpb�k�Q)+n��|�ʳ8�Y���H3m'�"�,��~��D���/�s*�S}d���A�����Z��|�����s��������3�B_@��5+wl�F�����Z9[K���q�� )��M�!����l!z�|BB�m�(w|q����n�#	5:4p\=C+jp���w�ښ�7�_�sx���w�#ђN���]Y?%�4������Lsiz�m���W������u#\��A:)|� %m��7�|��ZEq���뤷>�#�5���pB\69J��KHDD������\��5n�V�~�7��lUq�c���S};D��{�&�����������WAb��gT^ńz6��N�T���F���d;���k�#�ZBH��{��H�X-}�$��;�"��"���g��I�|/MG�k�N��u��߄<i��T_e��s�n�(`
�VA���R���v��p'������~.#�1_pydn.��Q{Y��D5�ZR�#�.Wt�+�*����I��SJ�'�E�f#���� ������t���Ia��W��Ӻe��|��dl;�=�Ѣ�����	tZ��?J����:��18������30d��;;�\�ݶG@�8�	e_4���QS;>
���諗�/B�BM������'��v�Hm(; ����j*]�׎؈*^GhN��!*���S9���n�ﰪ����B�_�f�f�`�;E�  ))��8+�;P����K��l�"�.�c곖vXHc��L{��St�Jxom���Esa#d�%Nf�_%�_�O�ȶV����뇒���'���׿�}L��@���e�+��+G�~��7����/�h\Bτ3o���dY�0�:�%����, ��{Y�n�v��S�d�FR9�ǫ�m��+v|�2=w���E�R����1��9�DAx�d����	�1�R�x�I���z���Ud ��N�.(���Ӑ6Lp�fs�[��9N(y�i^p��/l/���?���UꀒvI�MiN�{%� �DL;�{hHW�/�g�G�	��W~ϼ��u�N�q����1A�|�+��.�ײb
��a��B|Iy+wG�����mkS]<��W��(%��^�z�&o�������n3)�F���9Фx��W4�Y��J�^
�|B���-�rښ��0�����-���"D��3}1�O��� �:��1!���R����Q���vC�$�z�]_O���!���7<�AX��=#�:զ��j�B«�wK/~/�ܙ=��D���80m�S�9�0_�:��X+ .M���~�������he�?�%�ly��t8*�����U�����I�I��_���!��J�m���9�e�w��ش�E5af��W���!]5,�i��zbF<���ـ�	�s�7P�b��{��̑���>W��ȯ�1}|�[Uk9Å�s�
�ƃX#�{�"�����}�#��JTĊOo3'��	_����Y�u��һ���'�:����Û(�'�:��y-)���C��Ϧ:��LW�"XT9b��;�cϰ��F5�O�y���]c�yǛ����Г�o����ב�s�_d��f�s�U�P0������ci�8�-Y��$D�C`����1����ZsXQ�1������\1��'-���(`�A��E���X��7l'`N��l��r������^'e�Y�i���tx@?�R��E(����]�֌4��)���5v,��~J��k�]Nԑ��m7D�������b����)���h*˽W-'6��m�jk ��ex��5�j�tW����!���7��J�z�Ooo	��=B�\�֞���/���H~�G�o��v=��+����4�b\��O��iW���q�����It�l� �V����M�����q�l �~���y�&
��#1��|�p�?�0�d���*� 9��*���#���F�fB96�C4V��y���m��=�_��~��kկ?<��m�.[|��ʪ�$�F�-�?\_�=x�=Ц��'�l�xp:@&�qq��X����||�T�hF�!�w�=��g1���1|�;�I�����^2B�S#����[�T�ۤ'���	����|�;�є��Y�9<�:gE3��;�]8N~*�f�~�_�䫜Bc��$��.�5q�Q��9Gp��ə4��~6��)�S9qz6B!�{��[�	؄~u���Щ���GD�2%3z�{R��<��w���|�F�[(��S.�[����K��������?�?ޕ8K"?݌~T�m�x�oZ7#�];��굄�'��2�˚#5<����I��y��n����νY�M��'8�D���=fU��$�<��RLd������F���75&�l�J�1�1w
��M�b8�"'G��	�Ċ]���#k"�,������;*6�/��1,׮4���(���"������.�?j���Eq�����@��i?j�!ƒ2#~��i�0�����{�N�r�s��:�E����TGJH�x3�k
c��箔r_�s�ò�H���0Y�����$�:��V+����..F��_���SSO��&t|��!�׍��G�=�2�{��ưk'@�vv���Cpl�K3�	��_��O�6'a_n�pT�RB�e�j��Y��Um�9iT@�K_l�Ö6��� 렾)H�|�ú�&V@���P���-X����g�2f�Z �Z�s7�u�{s��،����Z־ID�����rK�ʊ�r#U�eҦ�~u㈛�g�I �#�M�l�Y������v*6v�G��q�|*<Z(�븋bu��r����sc�Qɍ1�4gފ��օ:���+ߕ�%��`3�+�7\���݀"L�,�X8@� CD��@0w+���K�6������	B7o�RP��3�/=�P��V?������6��o�k�LJ��T-o�v͊[v��%I"]���yg�՜uJy`K�;H��3Yc6¯���(m��w�����՞n��a���T�YS8�:��9hF+��u�]X{?F�H���O��4���F@�[}�
�@��s���7�f�~0��S�-���/�g��(���@i3����pv�iJ��ޗ_�H՞��"����ѭ����$��?u�ES�N�a&��~N��B#TH�٥�{Q^w(q���o^G�Tf-ҚF��B,�/��G�nc�@������g?���n%�\�/�-eO�j=����JY2��!���`�ej��� �+c{ <J�#"h��蠧�oͩ�'�YaTą�{�T�=q4��0!�d:V]���X�n�M���?�&Ng�qD�&$��H�G� zu5�'N��5y+��֍KC��v�O�[�;��
��z	��N�σ��h�w��`�%���[��v�]������ /+5O;�U�"3�C�G���I���n��
6b�kˡ��K2���v�Ip��b*��xB��=M[���%�CR�.���q�T)�,+�4�Yɍ����D��볯��C��&��B`ր���13wOz��KŔ���f��Zk>�x*���v���S��kmy�wӶ�}��8	v���=]ћ礨N��5��㤖��G�1�����7�&��%ٛ��V���(U�Hx�����Yq������R݀� ��F�>�وR�w���E�Sx��ŕ�U_^�;�7�tu�X����|�����F-��[	7U�����(�|�)P�zw�b�R1jB�1�J�7�OH��a�(����1�2�H�,o��Yﳢ�x֑q����0j*��)���
 �&F�)aA�l aO���ņ��)�1�����0�$����򓧁�ͯ��a�4bk+-LsK�b��(��w�U���^u�~��i�U%���93��2z����(5�hz�T����ٽ��&č��Є�ـ���e��)(3���J=�8�MH��	/z�l$�7HT5����,dp��v����}�G�Ay�X^��XX�_�Y�W���*?L����n�cm�+h�u���g��*�ډ0�k����$@Z��:�k�Wv��36�[��X�P�r��	E�v�	�O�^�|�#������ڤ�M���{R}�̻'m��ل�]�9D��MJ�D5��9���aY�#?E8�(d��}�ʖ�>����`ǈ�L�Q�[�:�Cs���\$��HZ΍��:�vJ�yM��Z�����4L�#LK���<��m_��7ω�		مJ���V�}�O�#��e�}�*��Z��ov-O|a����n3{���G�á�cn�l� �M�R���{(]�\:���R���c_ �7B����:���.�$_���%S�P�Ž�~�"�*@���i�Z�����ayts����h�s�,W|v����a�����+W�������;evVw@%x������FS�q��f�iqEX�X��Hx���M����ut�#�븦zHYC٧����AWN����cU�^/��pF��^΀�f��(�ss.���? �>3�{JF8< *�C�qj�G���,;<3�����-��֔��;�E��uyM�Qt3e,wr'~)�`	w�3�b{S�P��|�������ث��xL"������9؂-sB㇅H��C)�Y�j��Z��������m��[�f䇏G�/;Y=&��� ��"p���I�/D�W �j:y�#�i���3 ��ԓ?f��'B8������Es�M~��c� �6R���n��JI��[M�g��@��6/Oh2�=�8�6��K�w�{�>I���ҽACQ���{��]퍐�!��)��p��#���d�A�alU��3׌l^�SJx�[iH�G� \{�u̜��|�P�P�II��]A6��A3�{���,Z����*\����qk� Ĳ�_dhx��2Xeq�ւ�=�����L�c2Y���=�呿_����'��4��g(�������Z}6�C���|1ٜ��0`I]��V��c�;���/L����Ya�e|��"ɓ����uz�YL��+F��R�_r�?p�?�(�/�QC~���50��1�Wz��u����,Ï����=u�ox�b�	u�`u�8�0"��\�W�Ҋ�V��A�=rI��q�����o7���|9x�Ro�Û{�?Dז�P�E��*K��:�A_ţ^�����bT%�G/Q���s�&�-�.{���8�a�eL/�x�P��Bq����ͷ��l�����r��n�7#�=9 ���hS��ľ^�ޒ��S��*З�Z=�v��r�� 8���T
Y�xI��>�F)����luc�a��S��"=��J�s˩?Tw��A�w��Fc�;�t��*���"�/f5��&(P~� �V��r5���i�s�3_�C]��*M�v�(*n��j�S�4��9���g�����u��-B���,q�J!�g�F�S��噀�93��@�Y|`>�+	�CK	4��>4#դ��Wc������_�^-Y�6���"�e�m(7geŖɹ�YB���l?�8���B��m5����U�ُ@�����������6��&"��m�V�����c���M�фP��ó CS����z��nj�������
ꘕT�;�y�m�NT�=׊��� 6��C�9(ľ�zn���nn��t}���w�<�m�ǰ^j��m?f_�'�
�z� -�-�����|ˑ�r���D�IC�#R8~����tȵ]�/�&��z*�'{.���;��(���������a)i�<zVs'	R��}E!��9:�J�����T_v	T��I��x�*9���Ai�ʐr��	�oT���H?�wOOh�����D�#�[�'wvل�ߎ�Fg�Er�ᴈn�ZH��oy)���/�È/�g�?,�(bNAC�P��f�pS�&G����|<K���]a靿wKz?�L�8c��ݎ�������Q;Y`G��x��}��B��\�4�vs��V��u�qERhX �wz9C���9��@n�8��AН������fh���M�&�AF����v�4���{x�x�{F���J��l���X��̬����+@:�Ӣ�� ��j
)au�Sm����ETQh��L�T��������2֥����HF)#셍E�Q��䫱������d��w�TAA�M��zn����᧡��lw��RA[[���n���Д�yC���':�d5�C|�\���4"q��g��o�G@�0�#���@p���T�z�26Q�_�I���� |��:icl�:W��W�K)�b�1G���r����>�k�Z4��a��+b��&��ꋀ�#t��o�!56�y�V%�(w���N�{�E
�)-���;At��,σ�����w5�U2f�<x+��Zfv���ŷ���<��ؚ|џ�Y��=e��&͘{h-Gd����kiL,���z�r^:	h{�{ �T�L�	S���ŶM��V9E4ARG3��O�'�;^hV�=
��|�7"|�
}��u�����R�:|F�o��Xf�ҫ�@ x@�����d��(]��v�%-��k�\HI�8�JQ@|(փ�S��W��SZK�5\��F����2S�^�bݮPjUMx����hp�v{eM���i{�G�]���߽F�m]�0��{�hԯb���̌���Ӕ�g�C|���~���I66]�~�J:T��L��C�ױ�~��^�f�-�(%����?&~�a��Q1��tA�y{R+e�\���I�Q��Fz��/�8�3�_Lp8���b�W�Y���כ�;=��'���ے�`>��g/z{�3�Nz��IZf���vTlsuǄĈ`N���P�%cf� [ʀ�������op��qThȱބ)`+I�h�c�$��lh7���֭��EM����y=㼃�/���H�n����w�(@ؓ�!�>���&w!2���/�"��9_"�:B��
<8c��σ�i��[�Tg�����qW:�v�7$��;u%#۴j؝䵻��;Um=�Mق_98-�G�H�	��� `u����j���rU�X���Ng�P���3ٚ�~�梔*��n��G�֫W�o��vcY������+wމ͊��}q�Q�t̕���_�OEL4�:,�cyN��{%��s�	YO)�1#�r�uw��{M�[GdlV���T�]�˖���m��`*"�$�F>�xܕX�~�E+�0Dsۓ���E�W�|��ÍW'����j���B�>Hf?��)��c&���_���|��D��N���D-��_GE���YU�|EA���,~�ԓ<U�wx�����\B$y��_�\�f���-h��:F�C�R����mb�>�H�s�7EJ}��`������+���!�>�/̠�ѷ�7˲B�	y����oQ��'�->�\�g���2�Uχ[��2�8H��x�)��C�$�X�����x��\���75k���K��5Pt�/Z��	B�m~��\��*ɗ�+�Ryۈ��<E�������+G�(2e�NX��T:���Y��f�
�r]�Kb̨�k��p���V87�����X����q6���(�U�w�'�
�]���yqk���<v[>�a�ʂ�k�W��z��ğ��%y�נ�y-�HN�O��%�^�"���K|�����W�H}{�x*[]� f�r�x�
C�G��� B
��"r�_XXO��M�	I*��8�6]Lp+��'d"��b(�3.�j�冡*0�뵛��A�EP��E?��R�������ͭI��ҳ��X��^������:�����N�}�qӢ���ٳg�~�����$� �.�p���;3�~B�}¥wW��#�	��^\�/���`�_T����
��E������e�ǋ��R�S)���Ԁ�f���[K	��]��/R��߁Q�����0T�{ ������nJ}�k��4<\0��0>��F�xM����|^�>2�g�Ikrs<u3�5i��ҘߓW~^^n?O7�˺�'4�i!zR��y��g�x��F7=�yd��0{/��g\�;�u����2���z�e��ޙ��IU'�b��Xdq>n��I�Y2#KÉx5d��9]®������T��8+N$.`��>��ߚBo9���m�86��S� �L	#&�G����`������ ��bn���^,9�_��U��_�w���!�'�ԭ 	"�E�?�"�]�gv�E�V��*�;�x)�{3Y�����7	�0;Y��:�<� lM��WZ��=�j^mUb�t�x����w��dN�����֚7�|M���[<A�g�&���,qj��i��VS��lw*VTRƞg�$ދ�w&$�g�x�ܺU�����L29j�(8�>~�E��9K��ظ�>����t���כ��v�MG�?�֋c���=���I��'C��T��'���A�W��q�Ԭ4;�Y�n2����~��ht����v+�ݸ�Q��������~p�9��یv�^Yx�^�����L�p!��Oݾ�k�e7��ڟRJ���g�v����?�~�Ƶ9���ʛڙ�K�L|���I��H1���3�Ƨ��E)�v����K,\}@������ɉ�鹴86�AP�2Y�ՠ�\n���K�>U�v��><q�.a��+�g_)y~2���
竫t2Yj3m�sp��r�ٿ�S�R��?�v���h˫����-�\�ok���ߘ�O�i�k��*6_�坸�l�]?¤�*�DO�>����c;;Ox�~}�&iӈ���m6���q��P����l�
Y7�%k��U�P��d��#�X�6e�hQFc�[���R1��̈́���������{~�<8<�罿^��sfLY��������m�Rg�!Fn�"	׸�U��|�z1gda~�o��#��PQ�T`P�������r۟b$��ߒ�=��x\/J�� �� ���A;�6�bw+��zfJ�*�DE7�9�����:D��dޭ����_^��4����\��t���>j��� |u [׽oS">;��s��Ω饕[�h�4-�D����I ���6�n|�N�+n^�\����,���z��C��|���I�̍��{���f8�o�����Ȑ��!��Պ����9�Q�䄹��Yy	 Y%Y�"���7�<�|m:�<�z��U�Ǩ@�˛��G��ɰe�@�ac1Ǌo����ˈ۱�~R *�_w㹋�͎����O>�mJ�����W�JO�m������C0�[-��t�!.�0K���5� ����9�m	�A�J}:v�~�oh�HIS�T9�?j���/[�g�PL�8;[5w���PaEa�x&�0�r�W[���Ս����l��rO���pf�We�}����K%��e����yJL����!���j}y�X�o{@_*�;�կ>���ɇ偰�g�L��7�H���.�tI-��Y��9��+e�C�j$#7�#;��ך��p�������*�}M�|l�_��xK{�'� ��	\\C[����%��݈>Ǝb`�@c0����?��ZF��7ed�0��`���������l��~�� ?S3�GC�A��l ��)���xޤ��!AY�۫#�vw6�*t瞿�\N�����3ǔE�m��3{4)y��Y�Q��Y��/��:Y������(�c2��1�$�l�A�92����f�g��&K�ѻ�kD���|f=CCZ�G�y���+�B���e:���1pG�
o��W���g�;�����7�Z�ф�<�5�p����!�M���*�{3L`x��dCC{má��������� 0<5�K��ZaU��ސ�7K̾)5%�����=���,P1�P�f�a���r0z�-�@ �W�}�X:t�b�Suu��?��	�>��O{�+�(�K��T����M��]����6��@��9vYӐ�m�����$A ��t/c]N_pض��])n����W8������`%�6����=������d�����n]!�u)է콎P�������3���v�5��t��Q��Kb֦8z�}�׻@|'&�䶎ĶVJ1���g�sPuΦ�U�|~s��P@�x��z?�?/}��.���~"��c_4RP��� (�|q�p��Fk𥉟�_�0��ǭv�#�O4��,���N�B�E�W����h��uw�0:�^��Y�1��T0�[d��ŦM@
X��k�a��SU���"��@��%��tn�
������A���G#""�5fD�{��_��CdQ:������
��
� ���ӷwɖ��c���,��D�3����aW�C´^0�02�ӯ�%���ֈE����i�1�O���^�m֜1k6�5X���Q���FQI�2SE)2�$��/�I&�)�9��xE�%�ޤ�;ON��D�̡�(�Ib��%<b�M����������p�`�F�l�{���	���G}'�f��9�E�X�	<��ؖrIc�_���+���m�+S�y�z�sy2{�J��TnΩy�����i�����4��B�HX�$��=�"��g��r߿ �x�,�\Wc���$,���a�Ծ9o&�W�r�%S�/��#.M, ��o-��}�o��Ȑ��j�0��T����<�ҕz���b�(,�� >)j�
��
�}�3��n�L�o��Z��k�<ֺa3�H�fH�2%���Y&��f)P�.�*���DPf�;�wsU��#1��|�؝ۓQ� R&�Us*�7Frv@b��:���6��3"7���H�`k����m���$jƞ }�Έ���?�Z)����#y�iξ�r��}fa ��]elK�ue3c�}�b �]���P/�Ֆ�����Ҋ�{���%0�ii)���}��E��;��9�+W�meXX�z�>p�<b�:q�|q�%v�~%�5s��{���ƙ��[[�#���U�_2�����$���i�$�n~�~64'3�:a3�����M��ʕ���(Y��*9�!/V������_���
�⽕� \ON<�d�� 7��Y/8^�L�n��	�//=�"_ؕ̖��8�R'8��x�Z*=ݙs�_�F�> +G�N�-���N�.v�L�����d���ʓgOk�>���ie����A����?��[
�7����[Y��ٲ����{aN`�d�����)X��f�`�1���]G���'5�&+)�:62a��[o.=�:(xp�[v��^�5Ǡ�l��@�� ���V�����-JB?wn�?{�1�L'�{&:��� ���_�5�p|,D֥9��Ρ�T+�K�[U�|�����hS�"3���������R����B)�5D�#�m1BS��ȎB�������ooH��mX*pQ�N�'\)iϪcd���>ܓk�&X�Z��ַ���%��r�W�傫�~w(Q͜�W�CX�t__�|�Ubbf3��C�����76��T	fK�Ef�`;c�]��Y�e���'1�	��������aw),����})��ks����,"�+��fMg�I}�i1[��ck�`JZ2���1{N���9V�u�:Q&yH�'ih�7��������g���8M���(?,?�*X�0�Bp��4-y�U�ND���D��Ḳ�/nC{L��y�D>DF壆
�������?��em^޷v.�	\5��'S{��^ȓGPز��E:5&��4u³6��=c`����!��9��F�Q�@ "�H��!y��t#��I�=�>��ٵV�hˑ�Yf�{ն�Ͼ���e�?��rPpB-����r�x�3T~�����f,9���W#i�ELU��e4�<hX%?"�p���+/eoަ��BiȣWƋ9콁� �É͖<�ð��{76��2�����$r��ʯn���V���2Y��C�n�kAwj﷗������r\��=�����A�#�c�ж�P�Ơ�"R.����>��v�g�YT�k�2��b�M}me��4����-ibv0F�%������@x�WS���T��俑i��I���Aǎ6f�].;4����o��03���*Q�R�J.ua�G�Zp���lM��n�S�Є�/�Pw��|��;t��b��;"ȉz�9�r;�6�}2*���wS�p�G)'� �㬜xEڪ��݁ߩ��Ho�&T����"�ƭ�!�&f��b |('=��&���1�fZG?�)�,6ӝ`�Ek�J^����1>ah?���I�����Qn�[�䝢a�0�٧��"ߝ�x}8�rl���DW�=|-E�
��?FLhzs\�d I15C>UCڠ���$��F��j�� �:Ϸ|"��4�L�6�E���t]A���:���,.w�('�^D�'�
*R���	�8i��l����)B{�����)��%��9E#�SҠ?���5��Βnf�L�"\��jy�vi��D�H�}؃���x1��C^kZ)�)-�ٱ)T��qtp��I��i���(���Q�*����nAj��VZ��-���������;�l���	��V� �!��,>����pr�� �^˦�� �yY�)���!����@�{����y�0�P���]��g��D�b��/��/�7�g-�,�F�;#�1�����B4�ԙAv1�5*=ƶ�a���CTN��b″$��6��G{�|2N���f�I����TY���P��E?��{�=Q�@��q��O��{��֥h@�!�>��Eq�s��'eɈ��d��uW����)Zfd�/���V:tFEqZCǙ̡}�_m�%9���H����Y�6���N
"�:O��[|�����op�
�� 8p#��>zn�	q���,�����������u+���-�P�T1�M���i��������[_���lĈ���	��]B	��&LGRj�*ޓ5��r]�0Z60h�<WN�k;8�o�\��{%�擛���c���Y��	a֝:�(���烣P=]���5kky�.CO�3+��C~�`�ƃ�X����������	�2�x�!"nG����k]�!�$-=�� �Q�Jy�X�V*
Ol[�/��*�4�-tp#͔�%���@(-5�����ʎ3:�"CJ����䵛�bN�3�Q"�9�#��얇� �����4�3�fVX9�6x��䨣�Ȗ+���S�u&[�\��c�+��ii|�;���-E_%��4
��Q5��r���C�����c�28Jr�X]ѷ�̖���Ё��ax�
6(K{��
�KT���Щ�܃�����\�~���HwV��U�0�tt��""�É���:�9M@k�:��q��sj���_D�F��cF����ǘʹj� <{h�����7�" �q4r�[��������5p݅P��Ҡ����_�"��k�,�	h�t�P�=���C�"$Qr8u����0#Y.Z�x�]p������TY/=���|�"
H����?�=N���?�Y.��f4m�T-0�i����ᇼ�9"N#L�b�D�p?��t_?��6ϣ�K�����44JV$C������a�(�� ��/�cm�_�p˗�7���r�����Y�y[M
,�i�����{�Bo�;��d:_������9C�a��DIڣ�d2I�"㔁�Av��9�*G�i�i0*Ù���y��G�Eg]@� �t(1g���G��	m�P��n���K�nبP�:���Gi����DR�Knp�f���>��}`��1�H?�^����R�I=vB	�7V������@�
l	�O#��Q���A��O��=�����qi�����^S-�)�d��S1V78V��������T/�2�l��(�s��d�
5G�O_�rr��<K�iC���S����gi�ڵ����"�W+��� +����lt�#��
����;�����8&'�O�\v�B&[��hs�k��I9�;��op���e��GR��bxAjolث��↼I�^�Y:X�Х-�Y��'=����&�C���~��*����a�v��B�o�-0��L=E^c����"�C�$��I��r區��d'� Q?�)��n�v������8�<,���*��� @���KF73�+fv��y7����P���E׷�͑)��b�1�&����a�0B�FJ#�}ۨr�a�8� pX�����em�.���[#��e)?��MbGO�&|!܏q���m�M3l��i��O=U¢��`9�����
պ"2V�a��Ӿ�?�c��Lb%�&�3,`;8,�A�\1�Z1<��s�*��><bo���km���o9��7wEU�=B'�g�.6Yt?g�@�u�r��������~y����ʭR��bթ&�u�z�rR!�8@{��/C��n����|�Fs�v&��wƝ�/�H��N��U`Y�,_��%|�"o̝���D��z�y��Z P�\�^}�5���5�=Z�0��S*���',�A��z51U|]��O��,��>W�<}U�j@h��l^�"���l��Z����U��M�k���B�.&:4�_�м#\%���곘N3�������T��]O�e���h�0h}�;���H���'@���{��\�-�������~o�t!Z"�����kM�n}[�a�����c�䓷�$@����f��BX�,�/߯��r)����u�h�E��6�ԿڡD�|t=�AOx��*Kt�ٲ�T$ԯ���r;���a�V�{���J��kx�9�}�	��^���8���c���7�����]���IO3�@��e�M��+N���PK   8f�X���  �  /   images/5d57974f-fced-4f10-a93b-7d150e366d9f.png��ePN��)�
�J!��"-<�;��
���-����P
�)�ZH���^�yy�y?<����ٛ�ٽ�۽�E����```+�Kk<i�')�>�~$�:O
�I^�����+Ϻ��4���dt�4-�<�]�1<==�Y;غ�;��st��9��``І(HKhy��y'�n������z5@���I*��},4"H��=[�俜��dVM��������z,�����L�	����S����q[pp�_Et�fe���9���y�я--�V�X.V.�]�����Oq �AA����;���%f0w���j����GǇ��E��0�?���RY�u8� ׫1�MMi����������X���M"���
8��:�����w(OQQ^Nz���V��N�A}}}�y��A_!m0����E� �����%e���#��CB{4R��/��}F�
�f}� ��%5EE�����=q�P�E��W">�ĵs�D���iuuu�����OGk�
��D�����Y���&lW���s��>ͬYŁ0V�/��"��I��	{�'�
���H(���o*�^�I�q�QQQ�s\U�I<����
S#�5c�7A�����ϯ$'���;�B��>��5�ׇRA����&�~@����2c���R��6=Z$�"�y��A�r�����^�߉��IJ	*�0	ua��JХt ��/ő8�1�4B�M����l30l&�^�w�ϝ��19�٫��!!!��c(&fg��2\��f`
�llE%%�Ǔ�Xw��1�������?jyB��Ow??1=������I8\���+ɸ6�_����9b��)�:	i�
�\F�c��e55�[�$�� ��O���Դ�����MM����q%E�B���!�Q&���<|��ں��(��輄.��ʪ��e�[~Қ����Q�;��*���B�Fe�����ܓ��[.?2��i�ج��3㹵��Ժ����%���ե��xbA�ֆ�)�js4�������D3�&S�p82R�;���w����6��C{`ek;6)P�![�%�а�i�������9����_�5A�DIu-����wpI�@��2+a�����h�l���a�%�\� �G俵^%ooo�R��Ut�%����)1L�Ǡ����� �=z��G+�Y%��t����T�hSJj`�����}�v���&�o������b��y1�r)p�/�T"�l�7]�B�������(Tl���E����!50��H���|R�-�8�����`9%e'�l��s�����C���� ���=��Do��K��M��+���J����`C9W`��כ9���7�{�K����t^���3=[QV������rۜ��%	~��}�q�b�SJg�]p x��L���l�BTש�I�'z�>����Ӓ0�]��'��A��z}R.vG��Y��<56�6�������Q�R��*+��#sgý���?�D��J�����v����2�~8�fȟ��J�^�Oє�~a�Iǰ�s�^[��kfs�<y�T�C5!K�'˽�Mv���%ǷH���q#�pۭ愅�#ua��O�n� �ډ�����N H�����i�QD����6���h]�<����¤��w�zv�"�n�}��X��o$�DI1�muZ	�#��b����sC��*�gcs�a>	c �a�ɤU��YH���[u�p#yP��q�sr����*��w��k���24�@^
%?̕�dX�����!E���8z���:�d.�TS��%�M29U��֐�AM(���(3E%p�W�2��V&v�[0X� ��m���[� Oێ� �����������!���X+^?~�BI��01Sxt��s����G�:�;/̉K�p����f�_��	����>���:Щ�+1�-+�2	Lq��@�aD8� ���P[B��l���h��R�)|c���<�����B�l�bˊ���(���_�e=��bE>�L��B�%e�`���
y}�Mb>�+H6̠J�u��ZE����/c�+f�l�a�#��g�~d2��
�hl¢����ɐP[��43�K����A�~��)�^$�~0���oss߈AҐ�k0+����j��S��W|�V����Y�$�/�g�!���E��0&2�������+�"k�6yZ	��ѫ������_?��'K��:^��~C��;e��J�D��|��Z&�]���(l�@;��Ӧ����t���/�.�\·p�@VϫD-��?���n���vHb`v��X��'�,[���|�U|�Ö-;~&���N���p�g?q(?��=H�YP��f���Eka������yF�.�_.��N�E�o��:�`�T";Ló�w	�}�5��k��F��x��hz�ߝY�7D_��{u`4EMJ%d���eXEepbz��Ds\����
�oJ�=BG�~�AA���=���l�ծ��?J� �;���B�T���<���G���8����ma�R��B my�-�J������U�Z��[\�f���Y|e?��_�F�U�H�o���oz�+j�����WX9���%�:	��$#�A��))~��dϢp�����5��/d�C��P*�:�}��oV���sL�Nc�VWèf�%Dom��7�E��E�˾�9ZG�Ӹ[�_;KQB���$�O:�9Y�<�W���S�o�3�P�<��iSuG�O\�(o/�c����-�;T%W md1MU�⾚L��%p��g:h΢uXcI��o&���O$�.D��t�2*�:��/P��x �CJV�N#���F���y�mb�r�x����3v����W}W0~�#��<�Wi4��P��ǳ2$�"ĝ"4�������\(�������ҝ���A ���ښ��%+�3!4��Q:�ۉ�-`�S���G�k���A �^����n�R�����ܘl�װ����S��2�W�\�+g�\��ɾ�I�� .���l:^����C�f�EE�|=�ϫP��.ϴ����bɝ�:} ������{ggK&�&�h��n������4�(	N����+%���%���i��7ۙ�RL��	�1�w����-����Kf#ǟ�'�i��J����K�iǓ��\� ��ծ���l({_�1ss}����!:>�9.ڕ�A��~�����\4xd]�DIS��ڙm���'P�\�T[��6�z��o{�J���u���P{���Mv;ԫ�F9N�6�$�#���J�DI�������y!!K?��/e�픥��°P�5�t:�P9Om{���@,��������)�D��·�oiچ�-B�Hk�g�{QPHTfn���4\6N�;"�����ʚ��cTy�Em�t�q{h,��f ���lllB�q���C�PV�Y��X䃄��3P���׉LbiŠ�C�߈]u$��CE���K��S<�ZҨ���X9��q��Դ*��>�
ƜK�ΡU����4�Cv*���U����M +��BQ(�y�&a�t�UC���#���P#3�$�D��)q�H��$"����<��
D;6;�A��af�Uм��ikC�b"@��5�Z�g�	���)�Ǔ%۞Ue��@��e~p��K~�ߛ��L�-�s�x�d4Bű�K�_?�F.=kwK�2��Hn_�*q���O��K�o�������I�ef�|�&���|���x6�U���n�Y��A��xK��g᪩Y�%�TՒ��qi5R�^����aMYރR.#���v�~}�?~�����Z���)Zp�BQ�,�~qY�#�W���^;^���t�L��0�Ȋ��ddVQSYv��<�xN�*o�y"�)���`�;3'��g����2�*vJȨ�^`��O<��p���f<��05� �d���=m��3�a�Q?=�̈́7G�&�J 7hv(�@V������Щ|ѦYQ�[�d�.��X.ޣ4ە��$#������I�d��!0���kqQ��C��M����#gzb9R^:�R�f\���u_@;/�MNKdlz����F?}���pe���<�D�t���O^��g���&AAYAu"{�9Ec��iRϲ�d/{�}ׄ
Ҹ�;���~�(%iC��:x�<Q��㿽�ɀ��i��>}��W$tB�W=��c�3i��f�n��>..nx _�5�/M�b�3�3�ua3Sg~z�z����]A�~g@�W��.O�QBHHV��w�4/x�R�;Ҽ���G�x}33��X��Z�89��Z���͝oy,�x}FٟH��A�?к6�:܈�3�P�r��O-@��ݞ�F~*��8�*��#$<VXcQjٰ��L�Rz��Z>�����d�W0{�|V�uw}�x���:�M�A��A�O�s��P�U���p��S�a9j;��w����O����<�B i����\�ʥ����ˊ���v�q���Ӊ�!L���M��R��A��Pz$.�D���������Kψ�߀yO_Q����K��M%���z�+���<L�^�]�����<Ԗ�Xo�����ǩ�C!$D��Th1�Zڅ�@������2���qc�Õv�tܒC�Q	�[�g�q���Ka������7S�r�h��vm�#b�7ם�q��ؤ�O9�Z���P+����>�/v���.Q�!��9
�<��FM�0�l�Q��LҀ�h��˝��D�)�fw����DQR7+On�ri%)�3�a�Œ�<���̮ʏo~�R�1�6}5FBdI@�(ݛ1��L�G�q����N�A}]H��Z!R2'�o�1�v.���.zw�͢BP�9
�|��"F��o>�W';K��1֎_��9 �32�,r�i$�W��1�_I�9���>z.�NZ��ml\�۞C�ט[�{^�5g���ʙ����WNm3爛�����'����A�c�2&�q�������KM���f,K{b��u5f�f;(v�C��1~9L��\�-ӟ@��`��%�,Rx�u�l�#1.^Y�"^�?E��v��m�����������)�F�NS�����E�A�0�8r
?|yn%m u���W���t<���>����)���ݴN1GQd(�{������@`V�e��� ���EhXx���pR%�`3p��R4���u�M�ƌ���f1N�_���n9T�����"ǡ�|�~m���w�Y����.hvzA�MhL�[�W+:�~�^���ť��K�`6�sLL�ū=�z~<!a!{�sL����+%���Z��F�mYU�{�jC��l=����<�gbP1�E�GI[�o�ER�ߒ,���*�e_L2�bi�t�I$��b��]olƼ�ju��T�t�L�~UGo\}Y�oъ�6_����gU����=��A��}H�־���F�&���i�ݯ�&��(tiH�d�X�U�!H�ТR4t��mi���ܠ� 9�u~;���\���n��t�{���	Ҫ�k����R�#�
��y�q�b-�3��e"��o�:��es�_�� ݍ�:&�Y�>�a��wB�ls�����
V��?�e n��L�L˛2o1}�F��J_��[�''<���pYOffЛ�j�G�u,�� .�����NnYV�5�w��	�'FV�d�$X޲�nV֔���`jֲW��\J��X��tE��hh�3P�m�N
�A-?X���nܳ�R��?U^�WU�m2.���S
&���"����{>j���;QP�|��F�����2>�E���M��v��
�ohؽ�99\ S0��q�1�*�m䕞��}�?*/��.�]=6����#A��%�V���v��ư�J၃��>tJ��9[S��=���)S"���a	J�o��!�)�If�Z��9z��@Sg7���Dfڀ����������ť�=�"KX]-�ȑ<��Z�N�p>��7�y�l)��/��|����?�}a��Ŵ����[ ���"��E)hOVm�`z#�RVq9wpaط�+�Y��*}��� �=���&)�i�J�P�����+��~]�eܤQ��t�wxx8� ��-�L�[Y7W�<�q���G��kN�QR��cc�Z�Ϯ�}�Ĵ�f]؂֡��7�FP��9�GyW�ŬmYa�V���Accrw���~�S����c�[��PX�����Zg=$�\�ʦ��^�h�w�t5��hS}�T�1H�@ ��4v�RQQ�p-�<�D�_�1&�C^Tf��{���jX�x*sߺF-����n��9e��i��/s���
p1���c
E�>���5G۰��R��,��w������8���������!R��P��R��N���W�T&�j lx���&�* 3��B%�&r�����7+�Q���xev�;��+��w���k��c��G�u|�\�2�6��á�c�Z�QKCS�s�ݴ��;7�#�"7��1����v���.À���Z��y4<�/��>��l=!�n-E�ǒs�
��Ε�INN��*�[����v}��kuu�t�zO�,	������𜆻�0�8KJ�����1�g�w�;/���~�s�\L`��
rx�U�7�Z'�'_1����B��ll��nF�g�'Q�`)�4'E�5*r	�Ͻ�m�倵�*���~E�	{v��F��:�W��!����^�V�۝����KD�\ӽ�C�������;	b�;�e��"����L�C\z�c*Zhä����y�zm-�u�]�<�	�[�H��5��_�D״,��	�w����kˡԡ�]���ᇼ�_2ٯt�5�E@�0c~���_1�%��,l�̮�'�����h�)E�i������뚺�]^K�)��zHG�>'�7o(+m��R� �8hI��Oz!�0�������,��b�7��&�Ҋ�,�އ�<[��+rj�%o��<V��q`�g`_tT�׃z��U��wU�{2i�����啷� ������C�I������C�Lg�Q������S���S9�_'�Q��*W-�����|�\��`�A _���� �*]-i� PK   tb�X ���s� �� /   images/5d7124d6-db61-4e16-b8be-eda918c3976e.png��csfMۅ�ؚL�m��Ęضm'WlOl۶��m�zs?������zwUW��{�u�3\^N   HJ�(  �  h64����|Y�� c'��  ���$Q#�  __�"��n��0��j�d�9��ʁ�F��V�#u7�5�ƣn��50��n�?�cm$�?���.��=~����t��&a�̀����3x��e#d���I��H��+j��ʼ�W���\������U�|Y����1J���0j<K��=���&�9�7����<��K�QA��-B!�[d��p�+e�c�n����뀿��T��!?d�� *8�[����_q?��LPW��'���Yx�w`W��X��ꈴw~��E��m6�Q��V�ņ�Wߌ�m����x(≥��\�Q3����ʻ�ӌ��f�p	v�AU�rn���ŷ�%�1�)���'��%a�sO��U���rӶӹ�p��"��w�ʽױ�{xj�㋼4�(��4���n��c�7eu�P�K��p���hv��{�Z�����q'���20}�_gk�3�F'9_����.*[G�6��j)IH9�X|nR�:�?��0!�@��G���B��i��M�R '	3���Elh�X]	�qӢ�����+����&jqy(>��=���������Ų�1"�����1�~��%�]0���N5>,�Oǩ�K�\���`n �2���P����b��m��[8��X�3��f&8����4]���UH<��xa+������0Ӈ�5e�e�B��Is��>�����AT���W�mK\��}=C��ie�)�>��ee+aM|�i�K=`���OrƵ���O>*$:9ݭ8����)!l��g�S`�:U��j�,�균����o/<KNj܊�}����t��� x[�nɤ�Zr�[a�}{�b�q'(��W���O0z�n�0��� ����tᗵ�B��
4ɑx\�^9"��:}�_��IH:)��۽B�{o:sN��u��XZ:o<��4����׾��I�0�M0���B|�k�y���0��p�<����X?|�g��T����&��9k��}�lb�F����d�t��2�;T��v��C���`U�:�8w[-#O%>��N![��}5O)�e۪�-'f��4*=���ƺ�~O<���X�����(�1T 4p͏���2v�*�icd�x�S�����U���|��k��z���K,�Z�4����q���_�Jqk�������6=��c��{�
=\D�fƃ��p;�u���e<D�$���7��\E� U�6�ll��-l{Y���DG���ц���@�Q�%�o��z�hNOd OlVw\��W*��B��NF�A�~��qv��h�����ĺ�px��L}n^r�>��RC.�֏���l>|�!lZsI?J�rn2||s�jlo:?j|� ��g��2%_��v�|li$(�7�J�\�6���6��z��~�|��n�9��W{_X�J��9����;k����,�Y꼚i�;�؈����s�&5�O��=��L)2dx��ϑv�Kk��+�>!��d��W��?r+����
��L`gQa:a�� SYֵ����b&m�D�0L���V'\D� 7�T|T
����J/����%�'v�xڅQ�G�I��d�"]����}4��}�c�}��X�Ք��(��]�E^�D]��f�V�|a�충g�#��^��F��m�mg��1����Y�G�����}���ږ������˴�'�c7��c�9Ρ��H�����^ T�q�����
�h}�݄ł�j�ȅ�TiT`M�U��&Z��r�;e�1�*��{�^@j�#% �ψ'�$wcT�l�)9,߻��L�'�"i�K�D �Om��ǝ�j�l���r��`��[ru˰|���g����\�Q�y��cQ*
�3�_��V}u�Y������-"��4���������J�h4bb�r������f�-S��e��&�46hW<��u_g�����M!�E5�c)�T�t����NOx.��1�YL��������܂�� ��V(0�6F�
�K�n�Ov/�X�cPCP�rrb�u���[��l����1H;nE?#a��s��*��������q��ULQ-s'������y����rСsr>�B#�uUK��i�}~ֈ�?N�B��πgN�u?dd-"�%���̥��[A6%W	C�	�����Cm�	�/��Ⓨ�Z���5v��#��9�v�7_��&0�i�2b�bNP1��M<`�v%��>�!4~��9|�'�n�p?���T�$k�~�/�Q�L��v���G�� �VK�����e��*�c�S&ډf�Q�F���.��iZ	[������+#���Fn7���|����.��w�^7��ziM@-G�W=�'���D�?�& ,�uMu	�q�v��>}L�|���6\�>z�|��=�Z��݊�����n�?w������m���3�Uv��)3\	���t�՞��Ѥ���d��N$!#��TvO�9�JP����F��E�G��w��V >�!7����y&п똌Ҝ� 1u�v���EDm]qL2Z����揾���3|V�U�m�Ax�ɡZ�<�%�<�R��d۾�b�p���W����*[�4u�S@����Ll;!"H;/��.d���b m���ֽ-*؋��W|9<�cL���A����H�p�v��Qkc��[�t�����4a�n�_.�6k4Ń�6NZ�����w�Ӏ�j�I*��]YD�G ܓȗ�	LO3Z13i�oJA��-�����MX~?7b�aW�u��i:���.��<ls���U����y4���'���B�vy�n��������7�P�bP�3W�}�[�K�-
3G��z�Q���V=��|56-Ż5:�I%D����1�I��Oc;���4����!Մ��a��XBWW��(ˠ�I|�siq��gkcc\KK�R5avV�T����i1B�T�PЎ�Bs���z��ζ����Tp� ��J�|�PK��J�gX1��h'V͞A+	t�u���W�k�ழ~����I�,��%K5��ړ�F�+���U�+���\{٧Y��p�O�����	�F{5⎊sv�gG���э�&�~7���|5zle�k�g$M(�{J��YRu�	F0�d��`5�*n-�.��:]�dY�K�X�`�U�?�B�E�����<��yV�h�U���X���XM�e��dI��rz�����O<$�rjk!���Wi0�1@cu�]*+t�u�x�d8?���؁�Mõ�z�U��w��{1�t�]�؀vC�o���kʒޖY��ԓKOSk��[떸�ʴ�M��$�PH�B��SI��/�<?�޲��w�ƀ����6[�_U�]qk8	���P�wq��k�[��½�Sv7z�Ǟҍ��q��Qp��$���g�d����Y��3u��鱦�4�T��gDY�����nL��cy�Ƥi�C�U��]���2r���1TeeM���G�pz�^i�%o����3ꅣ
��@"�|L�W���E�Q'�f�N����81qpp�}�=u�Y�>�����gq��w]u�d�v�z~}~xs�O�0vi�S��vd�/��xv>mjv��|O[7�̪�!��wE1f�Ē����ڱ<�����*
��+�A�sA�յ����R��Q8��d3!���s?�21"FE,���1����H��FbV�+T�~5��(�^Ey���ў�33B�Js��Єܿ5lR����gw�;N�A�$M0<x���
��4-��Q����Kͦ�ߝ+U���&�m���&R� 3�Ӕ�2�-�.�����W��f���$�"Y������"��݁� =�;��I>�}(F ~�!+$$�c���ʴ�j���u��q��j�p(,//�,oM����oʖ����ߌK��lq�!��"U8��E�C�n�~�B�i,5�z�C��X��m�^��럣`LP���_�%�/��9|ԡ:�v�U�?8qp��BkW���\��e�����>n[Z��5'��S����Ҥ[����.���rqݴ��S��m�?�N�Z-V��:��5`ٓ/�,oA��4���wƨVW:U4����cFk�"ۏ�C1n��y��e�h��Y����t���hs��OEL�����ZRjA)��cӰ�����~�uf$}�[8�T�m��P��>9?g���I {؅F��dm�a�c�4�N[���+�%�|dB��L� �͑u�9f�֝�����Vtr��ӓϣ��4ԁ���o����i)�U��3��*�Z�z�3����U�dǴ	9>4d9֑?�o�L%�ڎ(Z���ɺ����W,�\��Έ�_L��g��/��4�&_�7��ӌ�܀�β�@�a7#+������5�9���7\]]�{���:��|�u���|?_�����^��d֢m�kvޖ�]7���{�|j��<Jx���Q�q�^&���XV�RљH'�)IOCԣm�GdQwE����4�Х`���l�5���s?��2�q��$��w~���5��Xż)~��m�!u8��/$�TFu�qx�o �3�U*D1�jPf�#��Q�"K�<u�߀�q�� �>̮�;�c�u���B�.�4-S�萍
'���ς�c�qvj�vm�aw=��Udnԓ�̈́3)c�D��ڛ�xa�Yq�ŷ��,��n�>u��2ʸ5;IL4�L4�j�9�(-�x^X�l�w�LFDMO���e��&d�6���,�����}J�G�>t�:0jy<���iW��^��pMN�}D�5��S��6r��s�;:�����3i���k#CˉM=��2j�����	��Efv�j�<鸍�O����wX�V/�z��X� �� ʹ��Ҟ�S;�l�.CG^~�m!J�O�V�^��!z���&���H �u�Oz��Z��o�����0�^$�#)�:A�;$����Y��0���8�r��<)���iM�r�S���Ӥ��2}��.x��������
��K�e?���'��Ξ}83^��xz�mga�vj?�F �i�m���o\li+�}�a��^?q�c�uы��>��c| زj��=a<c��T�[���e#1�O���V�X�75gP��b���� �8=;�T	C����f`��;E�S��.�����r.�2N_�6�_�C�_�
�`!}������xR��H�ӂL��gT�b��>.�h���{b�Z��&R1�t�|lso� �?��>��C7*Z�O�p�	.G����a���#L�F��Go˚�:�Y(s�kxXvx]���]����ܦ�!Y~|���{�Xk�YF<�V-�J�*ǉ%&6�i��������mN�'ot�?��5�т��Ƈ��,�^�^�����ٔcImQ�Ah���Qm��0'������Lo!����E����/E}��v�z52%��RS~���g���"G/�j<*<�L#.��䤓���䝴{mja��o�O�n�l5�,ЛB˰�@\i0O��I������h�c x��)��$��\����?���I�vqro�C8�Ä�c�Nf�\��TS�|e�UC��.7�|+|�5
���3E�5�H�I%�"9�N2�j6�zX�lZ}�<�j2m�S�F�����6��'����uT���I�ک�ge��(��1lC��M#C��JN���e�f�_�OJ&���{�韔�Ih���Vc�y��i�ꔀ����I��J=���n�]���ݮ��g�6�Qna}��k��<&����s�د�h�@�Ql���ʼj�9ʍ;I����z;�K�r��F'���;V��,�#�����2��ˎ� �CiA�6D)؟f��FZ���	��'�V����q��\\a�E�9�&T8�_j&�B�����6�^����Q%s�-����e�F�ލH�G���O}�9U3��c���-��չ��`2�<d^�F �L�j���*U>��Y9��� ;�l�8~p�-�^o����F>~3���|8%ι��WW��ҫX�t���%� M��!���J�AZ�(�����0�_sCݩ#��T.QȦ f?�OcUA���Hw+�ι�W����*M��Ad�K���jH~+�aQ�G9f���!��N����D�`���e�Y��|��%�Q�d��
n�>\Y
�J�AY|���]�п�U�_��G����m���kX,���!�{�����&_��@�$�Μ0l�њ��eSS�c�GN���.��!e�~���c�����:��{Q�"��G���V����w�M[���uk:������!�NV>O!k��O�4B)�?���߲?����%�@Jg�����fU�62��(QT�\;�r%���MЉ�P�28[(���-P��S�;����Ȩ��L}i�Y^S�	Ɔ�J$[I�V����+1`�^|� ���L�Lؤ󹬓ެ�	W�?c��g�Oy��Zm¶Nߪ;��wB�BР�����/�Q?΃�J14�5h�~sA���X�
��e��Ƭ{�VT���9����\ƫ#�v�r����_�h�a�7���i�J�ƎE���FU�-�L)�9�
k/�Ǫ�.>�U{�y�� �ޞ� �o>$�����d����P��5K�1g��2ef ��NjE=�
.�5�MIi��ۃ������)��{�CM$;d�}r�@�w���xi�ʂY3�A����@*�#E�"W�&�b5�y��D�f|R�>m��I*{�b\<�]U�*%�VR��bV�g��_x�]k�"�@���@5�� U�q6!+�%	ۧ/,=�D�|�%���z\!_'^4Q�j�>�c%\(����.=�ǡ10�n[ˁss�Oo+�X��f�$hƤ�������U��5��|��M�V7ý�	�p#R?�ߕ���t'!i���p
���u�?G��S���j��S�B�q�zd@�����f[��a�HQb���_C3��'2�����+X���ze�����'$XiK���ďf�a��z-��}&]��ύ��P���~Wb��̓�hT�q�J7#�?'ޒ�'U�x�4lپ�$ʁZ0���<{1Z�z�s~p/o�z���NL!��6��q�\����E�����2 �n|3\d��d��O&��]|�A��Iqο�b��^�u<���"��?f+�h�c0�=Z��]B������9��ٱɎͶ�h�\k�*��?��Kg]~<��w��-�p��~�郘�C���.mêyq'��� �矒~-��<7��#q0���I���*]�a2�����$����T�M��Ha�H}��Ր�WjvL���p15�Ux
���&M~G�칇��Q�(]Q��I(�˴�_y}�[.7�]�D��|�,'�� ��+�}? ���S��=��n��|�L������s4��)�**�����7����ͤvv�����8��f�.��gF�%Nh�,<뤠�%H�J�rH�$d�
�V}��M�+gn����ϣe�ӇW�C�� ��[c���	x'��)�˨\i�հ�=���!M$I.iI���qu��͢����:?B�ͫ�����nt� �ԟ<)��֓�	��(~��.ڿ�^���|ޒL�tmJ��xz�� ^E�� ����zez3!�Sgu�¦4J��Uc��y������cvF��/�_�o|O�kF����)���;��m+9R�I^�Y�Ύ�����~��Q勧�6m'EH����0ޗ���%ن gJ?����<��|���oN2�׭1���cSΥ>fAU�Ϝ��->K�Җ�l��s�~����4�zc�]����o����5������6�Nwqc��a����6�f.P o�E���v�K����{�f�`���*�ϣ7e����Dg��t�]Z�x����ChY�gc�ᶝg��	P+H��p�d�0_��f�ع�k-�H�oŗ_�_�:ʨ���]]��c
Ά���̭d�K�̂(����W�I�d	��*-���W�M¸�޳{�ۊ�3M4j�y
����y�.���\��l��k�i�W�����A��q�BAh芓���.�fq࠰�5�^���0>�F=��5��W���{���ش"s�$*�τ�"�����T�����d8��!������:kW���}��y����ޟ�2�� ,�Ap�[iu4��G`�h�pɨӮ1(!��ф���(�e[��Jx:�H9��Z�U�on����Q��u#O�Y5}���Y�������O|���\xi�2�V�/m�sFg��J��0�8�x(ݾ˶�O��Z�2�oD⽟y��~\Q�}[]�<ݸ�y�8��$���NH?$l���P|�7��U19p���=��)�R��O.��Æ���)��:U���:̨N�g���s��w��!P�o[&Z�Y	V6� �uT6�ϖ�/�p�h"�D�b�q�6t|0ZoG�)H���@�6M�x5eUM�q~X�IrC�J&^���D'w<#q�KZ���1_�ԚMV��{C�3hH��Zޞ�t�>�l�&�x]7ݏL+@@-ɸәt���o���>����O8��PI�B�'	�l~�[ƛ�;6��L�1�,�'y�A�?w)�"���I˟ڑ����f���+Ձރܷ֝}�Ib{u���?��2{��"��7�|�uӡ/B��7������j�z�0����t���9��-�q�}�������i�L��t^^�?���r��zA�7�����&�{����A�RU�nTU%�h����Ϻ�£�Y��̆x{��_R�:!�}\��^�m�ao���ČM��v��<:������i�"�p��	�a��}��`���o�E$�$�T�r=�@�T[Od�ݴ�p/z�����:�1�roMR;Hj8&*���>�/ѹ�`�>��s�X������l����r�@Z�fռ�w9��铮�E=ѥ=�d��}��@U�F���W:5����#���t[���FJ��KKz�/V��}�T�҉PO[��	�A����9B��ղϩ0x�_0Sr����K��!��4Q�jeN���7U4�o��Y��p�a{=��X�AH����"����?�c�4�>�]90Be�͉S �/�-�x����v�eG��wm�f�w�%J4�⟭��Q$��k΍�P�r�CZ���c���L�m3�1�x��9��t��z/�V� �<�/E�3ly�c�F.�?8	b�}P+�B��M��J+R�
�4��6�=(����@�!%e��+ߴ��s��J@���DwIK��Z��0{Ja��[�,��迷��J�'Q��w��g3c�E�1������I+��ϳ%�7�\P��6q�K�ͫo$�R���^Pdi�*kPQ��l>&�c�CB�*�=���c^�J��5��P�\�
E|	����I�L��<��C$ ��!#�qQ+I�&J�C��4;:��,@��[�7"p+?����!�w{�w��<YV����Q[�@��r�	�Co�W�<�*y�ls�M͢�M%Va��
�~}�q��Љ``�7_}?�8h����'�C)�=R���&O�SۊϞ�	?��������2��2~L/ńT�Y�WΌ{�ɸ���eЉ�E\%q�BA���
,�/��3������K�C��*�fv!̛5r�!��D�/�#�QM�2QX��*3�۹���.����;���dP}_ߴ�M���=���@��_���s��}.�u�$MRdH��>A��ndn6���Q�.���)oF9�o8+���K�H2�Mށ/ވ��tL���ť4��W��q~Lf�E��-8i,�0c����
�2�y}� ��$h�d�Wa�����A��7�!9��jW��ڴ �S�g�L�;���05�{�-��X��#��b��+������ ��
�ԂYv@�q>!�3^�@�U�q(K�a��=�e�1r�&yGr��@�5�c6���p�(�
�ll�u�A��8١�[�?�ZA/6�>�5��Ť���f:E/p��RZ�bGe7���0
r���=~C*�-�^�`EH.񼹴T<��#,�"�p�R foR��a7ty�(�*���+Il�¹o�b��S��f�����l���0jا5��\�J�s2t��H�N�(�/�6�h'~�M��x�u�X�j��W���i7\D	h(�+Z5^����Q�rRE��:�p>q+����E\q��0f,��gG��9� &RP����I���p���{�(}�c�H��ˮ�-� P��H���*ж\";�;�[�(wb�S9�F谽"ݷ�A?�hx4��Ҵ���J~,tM�S����$�K
`�F�X�A���B���m��$M&��,�X��sa9!Ǽn�j		QL�ٓ����w��C2��);;;��{&=���2�﵋`�l�F��U�]�pI�!�f.6L�r'��'��Pۃ �%��)z�|"h`j���B5�����h�-�@����6#hF�G��ʄh�5��q�KL΢S2��1�U�Z�.Z��b����X/�2��a�i�M��^��8`��}Uk��Wg��jU#��#�P5k���p�+1�����h�oy5d珕Q��=��*�/��ZOȍ�wr�+�nD_w��-^C���X����r�ٓ�F���a�U���[^�d�0�E���k�n
�p�j�C���Z�Ժ_a�Z�4t��h6�8��6Yl��>7p�S*�p���G���k$3P&DݦT���z��]���Pe8�Z4�xF7�P'�h�`Zͦ�%�|�����T7���:�V�ˁ"%!  ��UHV 9X~���.����MGP$� ���0���B�b�U����8�)3�-��T�^��5j^\�$ݤC��d�T�v�s
I��`?a0�L��:�f�]�*U�j^��̼ ��㞚f�� �#�[��XE����O8Z.�Z��������!p5��+�%3.�Y���gn�����)�q�n��k>�x����/I�
����e�?����+���C-*�������~p~c?Z���
����-|,�Eü����X��7�v�`�t��6]�/��9V��f��܉�l���t�<T+��Ƌ��&Dɂ����ۋb�G�u�
�؎�hNy�:-->�r��9����װ��N�ςZ��	mJ|ޓ��DA~nmy�M�Mre�S[�o�#+���>���W�I�Y�p<������BK�={�cܯ��(��p��v��%0��c�-Ww��C�A�K��X����́�H���X�5ݤ8�<Hѭ��?]{�t���-�p��v�Ł��9��t�V�� �7�(���FlNFC�2�v�QQm�-�f&��ơ��"vJ�=O=�,�9{gx1igJ ���zƠ�)A7H����d��6�R8�����2b�D�
-�?��Q�3�~��&��g;�XΚ8~�a����(�8�Oc�7h��P�p �ˏ�.D`t9mV���V�� ����A�������F˃o6QՃ���	��t��@b�:~�~�CO�_���:Gz����Ď��������郣O���z��c�m��;��z[ ��n�@�B���sܔc���Y���s���JH^�Yy��l��!t���A���jh�j���JQ��vo��ISTR��_7�}�'g\Bu�y��
�fz�!ڪ�2�l1Tg%��wx �'�T�:  �K��'!�^��֌L���H-V�V�_�F�H	(fFtF����8e1D����6��#�&���<�ޥ/��.����X�-���m�l=�e->^n���i�v������f�_ h�����oAr�=�n��|^xK�J	�?XX<�aL�#�5`�(Ƿk��_��Oo�$���6� ��(� �Jź��U�YU�k=��<~�6I!�kvh=���ӥ\eDx$v���]o*/t����ol���.2���@��U�jm�d�!�ϛgվ�mk}���g���<�у ���q�v{�^#���[���3A���u�_|P��U7� (�m&A\J��5��u`+�..�^̕��S�Ӧg�%;*�4܍�:ձ��� Ȕ�8Kђk*ۿ�wD�bF����¼⠀1G/f��Ŵu
�6uU��)�^��+�+τH�5C������� �_l�4"�㸃�6�Q��V�	wqq�i݆�?];��{ +:t�ږJOo�t�ژ֞��>n3�_2^�zF���N@�U+��8��bV�*�A����d=�@�1��;�.̜��f�9Xd�{�*�:��H�Qg�	Az��6��%h@�?�.VB�$���C����1/I�S$�gf�=
Jr�y���ƞZC�n�\}��1ܓ�
��V�*]��m|V��i�.N�nTT��v�W��&@�ƙ��H� �U�P��Ȥ~�褠6O��km�P �Qm��گ����[�� �����l=ʆ�G�ձZe����b�%36��
u��N��{f,ʍxg$Jc+���+u�
Z�2�b�Z����Gǹ���7�)^ ���)�UG�,�_#V̧�5�ȴ
:U�]%DB�v@��`T��n���ǩM�u~�E���ώ!��ǰ���wؾ�@��{�8I����"�Σn�h��G{��8�O#X�,��&J�t��W�����y1�p	�Q�#��ːF?�6�9Ӈ��"�#D����8�Z�Q����]`��n�
/#f}0N����rب�h���R&�fP�$ ��T7��7[7|�:~�dl���)��T��_"�P�sVL|H	K��ٳzX&�0^���M��0�S_�ް櫧�D*��,��1�E���wj��̈́�>�e)<�I�@��B�����L6����wؑ+�љq	�
�2��mQ}/�7$��G�[0��^��~�kW�#�}8�� :�m� =$�߀>-�k�J!_S�#�h,���wh fL���1αx�lXG3������ҹRֹ�>�����u7G�E�e::���o���u���W/�����	��x���ۅыu�(M�TN��3E��q�qϾ��p��6\р���1�}H��*O_Z ��L�5�ڢ�\��ُy}zL��u�1��b�0�I�8;3��D��n��]}��~�7;HΔf���7�*�=U�W�]
����.���錸�d������g~FK��céը2͂�_Ũ��P߸
 (�!����0���>z�|���=��!�XC�k��f0^�ҳ�I�,���`�5�����[��C]�Ab7�L��'x�jYh�����-7�ӛ%r3�9[�!b�N8M�̫�ؒ���r�������i�Mv�.�Sa@z�!�Q*.V"�N���O�Ѩ��} >�gS�H�r>v�����IR�ӎp��q[W�J�R������UYNO�A+� %��eڱ�3@�1���W�Κ�����VJ��(-�����xD���U������ڃ��l��"N�Fb�_MՌ%v�줄fp9=ĺ��;ed9�l��X��}?!�:�p��0�HQ�� v^�K(e���ᇏ�������Ǎ-���x�96������T0�6v��a�&���j��a${�<�4ן��XK��8��+ȴ�܉4� ]�:��ѻ]���}D�z	[iIۂ���sYhUyY�|;fT�@*�Јѣ�օP�]t�M�'��u.(/\�E���A�/���7p�!�����Y�Z#�CM���ue$�b�X�63up=�b�i4��AY�5��|�9�p��6ēsj}6��z��U�,���;F���0Ǹ��C�9�����ioX�휯��E
˳ML�ï_0.�|�/�M�~���@�	��s��Kpd��"B_pk�j�=8" p�:-�$R�@oG@$�ʚ��U�q9��P�  ��~��hlr4do��R����0V��Q�넯��<�85��wl��`����Ɣ��.���7���s��%EG�ȵ�j�G-�><8��ǂ��ˀE��f�}Mx�}�  Yvj���l�t�4�㠸��}P�U�yk���W�G���E� ��y���Hn�׈����BZ���C�`"*���ϝ)iv�D��v(,]Vt�l�)�n�JQDjBwx��_���<�	#H�nWMQ�=w�}$�� ;�,mR����������w�Y<����,��1�*0J�J��H8P�Ը�Bc!�X�#Q�z�@�>}\�%zǟ�'&q&�t:P��q�*�7�ԠS�lV/3��-�%��.P�����C`��t&/4��i�8Q�P�u.e���u�l��q*8S��z�GY��F1�M���$�&�{�����׊~]�!��|��ou�DF�6�eд�����v��R�3{P�:R�����M;��#H���WXKW����x�1Jԉ< ��=���dm��C�2��U-�+����h=:��N��
'�LQ�/	�'-�~� s�ѣ�k��.�N������C-�����4ʞG+!�5گ��1E.�c�:*�"B��#%�4��=jQ��%�A��n�³�c��/������Xm�MPT�CD?Ȁ����A�k��ʑ���.1�"Q#�
�Y��[�.Ɩ�Ո@	�R��2D���R@9�Zy����F2�DA~�,$�6�c3��촟Z�~��
���d��ㄻ�M՛"�?�~�:�w�b"�x(�$�	������K $���7Zϴ�ynP5�.d�����9�E�0O6i<�����GB{s��cqft���:oa�+B&&��>EJ�A��9���p�,p*�0|��?�ƺ��G��04ɝ�nHG��
�ϐ�[<���Ź�I
�U�5D�k��e���!�����#0���f!P��h�U��K�xTo{����_�m���>Y��v��݉��w;U���Aw�Q����@�{@�@��V�[i��=������q�:�Y(FNM +�مq{+7��_��Q�<���-5?Pa��k�hdv����Q��k���|I��6�� ��TƟ���ؠJ����򹊩�@�L�`�������V�G��]"$�	7-lQ�{q?
ZUβm������רu=�PS�%qs5�?BA�մ$f@�Z�Bq☘4)�:)�sK�0ȝx٘�BY����"T�5#��bDe<�f���]�N� _��1�Ed��=�Τme]��ńV7�	�h�z?d_��t�}r}�~�4@�<�i�t�R7u�
�\��]�F��������P�p�a�1y�'	?���W<��ş�qb�H�~Њ+�#��tf����!�+6��8K�����5vG��L��|S���T,�f=��I|L��u��j.��U	&��5ƛĄ���K�][�L��&���p7$o\�Sc��̸��c�o�P��uy��=��4$i��>z�����^��Itv�6�}�ҿ��/ֿ����d��J�Kq�"K���������F��ݪ��$����2�{�q��~�2Q�=~s�o������ r[�ڥ]�q�X�oG���{e�XNn8M��uJ�?�tcyi�v�oO��¹�z���}��ٔ��V���i��0��i����OhE�b2�9����q<wM�d*J��"W�6L������~��AH���V��7d!S��=\]AlO�|ތ��V�-C~������v1tI�g���m�4,�I_*��DЩ��J>�<����v^�x��k;�a�`m��q�~JQ{/��YX�3�����.�d�)�w�y�m�Y�����n{;ץP/[`*�j�e�[dͬ��n߃�P�I�[��J9ل�"4^�Δ�V1a$~�y:�!tل^�+�G}O�����VBઊ1D��6�<��_�rImjα��Z�6�2���s��d����08�� ������Ao3�xv�g�{���R떩��k�H��<���Uc�*�[��G����mF���T���V��HǮ���]���X�Iۧk��,�D,�����2ӫG���x�f' �{���phRF�纎�V�����4ܣ>�����y�e�%~�h�#J�B��w��dd�$0m/����Q�:~d
|I�ꯘ-%��E(r;{�vϼʹUA�����v2�j�%�tdεrVD}�w\�P��m�O̲9��������+l��4O4����).A�O�ʨ2�d�V�����%���)��͔�@�a��W����V���т������O��J���C@���H�GF�ʰ_����X9�����/� ��,�ݲ�28�yڗ���ř�?���������DEsg��N�9M�Y�l&�VD��Cv�K.�Jl��
�Oei���gK���tS웞�I;���a����Qc��M��ҩ���厛&�
�as?�d���	Nd�N�vi�Y�0��A��J
�?\A'��������;26����;���p�tW�f
o�B&��Dɮ���](����J�-7�)�,]&o��*�Vk�o~Ov��+a �o��Q����*I���W�v+��&9xK% l�L@ �c}�E������N�6���L�a?�P���lU�dǵ�52+�΂p��s���s���f�463�,TX�d��;JA�7��:�y��S˪�eJ:�%e�xf~T�s�/�.7��!_L�b��J�1W��P��o}P����NUdd�!]��$T�����ؾ���[Cz�zd�hU��?}K��/�NB��%-���e3��dGcE<�K]բ��Xq�����
�����6_FY戮Vcx���,>eW�PWؿ���/٫�Vה~�7&ܶ��Y�����~}���v=[4љ��Qe�I����x!��%QU$zaO_ᢉN}�;��2��o�����Gb+N�ͬj�����hM*]�$|�T4��l���X5
r����
ul[!�wr��G�e3��9JqI�&/�@Ǎ��U�Pp��7�3���n��O�Oy�;A�2yb�ؙȚ��� 2��P+/
�L��j���6-����g�QR�����9l=��v o&;�.6�I.�����8��%OB5$��̸ה����s��&�D��bK��$S���ׅI�|�$9��gZ��T#�MC�]�TV;�s��L�2��&j���3�*��%+�
��{�9
�$R� e�p��6�m����,V&9I
,����A�Uw�i��3��Ǚ<�,��C��eoۼ����&����7������c[?l���;�Y���5�-�2�d�'H�z�Y8a�j�)�ЧE��4���(Y�/`p��L�/ۿ߰���|�f�̉�o�ެ���h�8n������*+��`��F
���
��k�S��̪.���O<�-�j4��틚�Bݵ�Z����������D��1�݊��ZU�Vz�)���3}ie̵����Gu�,V�g��:�5s`fE�B$4�^�7� ���<W�9

����?�X*�nAd�W4��l(Qb���Slv�\�G&����D�'�a��d>Ɋ	@���q���X"}��$�π��]#]�i�ifK��zC�jQ�j����/�}��:f�(������Ѱ���4��Fi���n�đzb�H�GN]�fu���~6^�=*�dql`m�N!���ѾS鄓��y��!jՆ��Y�tg�Ս���0�y1�H-g�da<�j�ڵK�0�}CdόH�C6
��8��e���l[�[��%�x���k�a%�7�R*�4�(VaO�x	*y�S#��Jʄ����d'��V�{��} ��%��zRcp ��K��fN~�nҏ�4yPRU#)�4��+�X�ȉ��u���� �v��e�H�i@@�ߋR)�h�a�(���,�T�� h��2��?L"g����y�)8�������� �"2�ae���?Fr0�Mg��:���@K_c�-���x���1�+���>�Y��x���a��R�<��(��>�r!I�������R�m۶i*K 1];�S�z`�A�8�#-!��3�A�I .΅�"hp4"�q��=;|�ˎ��0������~c�|�JAǂ{��+��_E�S���0��c:b�V��1SN>��|rKs%Բ�'A��ۅ��Gsa���u��$S��Q,c��(�o{ �ɺ���������.d�kR�J�&�* <�W֬]�+I�T�Y�e:�N��6Lą����49� �7�t���J;���I�6H2��x�
���l٢yG ���q�NpEf5`�ܑ���p��\ԈfYKm�93�p��Y	��[��V� �0���A�i,�<l�
��C�j�bH���D;ܘ:�h�ΔL��4�������������c�DQ��	q�r�~s�a�<��%�Mo�\آ�7r�,\��;��cTǅ�1��;'�oN��%>�N�dOl6S����8]KN�SsS]-)���i��?����SH"�#X"�Ѩ�#F놲|����4�Zo2.JW�����SU�Q�*�
(/ѿO�e���Zo����X���C������?�����,�d����N�����Brx 0���&�s�� �6lP����5XU�"bsu�	��Hb��T�qR7)QT2�pT<8��Wi�`��������Y�eX,bڡ�x�k_����.���j쏥������yC��]� �u��cB��P�z�pH^�j��?�fy�:y�O}Ɯ�,����D��G�AlݺE6�y�a�k�I;&���-n��<$���+�V��ɌVӕqN�Ľ��%*��W�xq¼�H��O~_��H�
�C���[eϋ(1�0��eX�[��+��qҭ \m�һd���i�݋�a�~l�TO��o�,U���~�µW�8V�� �}�k�����`mJ/�㔪P|�����Pc �.��'f0�0���Pc�҈��l�����0G]
���|��s���8�%?�D�
���ZY"q�h�0ox���V۲ap 0J]#y�\����Z�!�g��i�J�u+��f�������xg,1�אѡR*�Jo���3f@�W�W`:o�T���?W����]2<tD
�b��j�>��P���XW�f0P3?����f9n�9�d�n	��9X��K����s�>��7� _� H�նo�A3���yC|y����Γf貔���19|��3�ʥ���A�b��.��K.Q�
5�����Z����K�@LLw�xu�ʀQPa��ΦƤ�b;�(�3�_y�zl\�#S�� �h�'�ö׋��nh|�%	�	�7Ζl8[gB�da>�.t=hVN@ðq�/����P��-oy��p�z��䤑M�n�lT��E���n�]�xܑ/<CN[{�T�jR�c�2&=�>	¢�A��w���$g8����^��hr9�%��#��NH�qQft��.��Z��J�]��ǂ�<Os^pS}p¾]g���s���]ق��Aw�]�Y��5	#�T��_��������37](=}+e���%�sE��Di��D����*���7�Q���p�
��&�^�O�N&f�>q k�@�Ŵ  vu���0��ׅ���،�f|��ya��R�to81�
����v^0g;���1�`���K����R��
2b�ep����s}���	�~pTc@lc�Y��KSy2:,���o�CG�w\w�|��~P���Uw�-[P��S0��]m�!�/j`�����5�r�I��(@�����c���5'����QvfLD��ᩤ	�%��6��d��~>��d��Ȁe;�f�
	WW���b�D(�Ұ�;�U�����|�w�I^}�:�$n���:2��1B�';T����'� ��xF��o|C3�x���cB�L��+-���4�j3^���s�9G���.�/񼸨n�q%3љW.xիe�V���͢��Au ��2�=�VFZ=q�`�X*@O�

�y�# �����1��� �=�EB�C��&�r�3v�z�/ˮÆ�#׾��r�Ƴ�H�\�=�R�%����*�&�M7��?�>�cϑ��X�~!��Z�Ɯ���L�)�SK�|��3��ɖ�4�C����$66PR��(�hE��|*��'�#C��� ��������o���$\Q���B�%m�F�9X�|�f��gT�|vK"F}0� ���C���j�ꆁ�Z dۥUki���QË��0 j+ �m�]gc����0�#D��GG�sww�,�]jf?T.}	����&�B#��J�̐K6&����� U4uv��^`� o4�u�E)(��`QEóL	�aG�Ql�j�բ�9G]�
�ɞ���W�R(��q�v�0`s^YC>���F(�rA�"��Ss��2�R3$���F��o�'ʼ�� ���V�?��@��/��� I��]� \N�1*���֌����<E=�4�����_)Fz��PS�����N8r�5o��V����~����2��GU`�����) _���f׈㱁'�_i�L��k�E�8p>X�~�NJ4��ڌ4�m������zG@�~\r<m$���u��S�݆	�c��ƺ񼯶���C���vyp��1C�AXN��6=�e�#H�9n���`��=�Z <���F��$U���h���իW�c��_UU\x��rҼÚ3*'��4��1���m��ҩ>�^I��7�Y��̘�4OE��(�N_+�����^Q���,�*�d���:>��
⌗%S�5�A'�|4��+��B��?���`��ַ�>���W�E��:^ ,Vʬ����	3���������ň�^���o�G�Ŏ�B�2Ci��P�HB�CC�T�uȆP��#�^�3o������6"�p\g^,;`�c��g��n���m�Ш,�d�-f�p�GI�RW�}Ǖr��uf�#f�n$���<z9�!mCL.���%�񔵬BC[OOY�v��r�]�I�5�4&�=��i�3#`�
�&|V*�R5P����w�m��,�l4H���"�5l�>�� p�+b�R�����a�TI���+gd��{�n�u;Y7�0xtl�f�p�+�&�rF����l���0�lR�,�	І \�6��a	�G����+2�z-��5E�Y��=��i�z�5[^�.Eؾo�R�a)[�H,訙�r}o./s�mFiƒV$B.�J�,�l�X>�W!�����w�������a�:�I�/pF{���p��+u ߫��Zə���L��u�8�]��.�i{Eثvb�]�3��ZT�;n��av��f�d�t�޽gwa&r��s��!60c����KVb��	t>X�}��j��1z�3�ZSt9a�8�l0�x���L��k�&kVwK�ё�ډF���U��w�j v��\rɅv��h]B��a��H&���W�z�&9p�jƴ!l^��ƀk�*X@�c�Ft�}Y-dpI�� �|���U�7���M]/�����`a%�&��z`K�P�.��L��8�N^!6�0c�ho���%/�̉�����C�>�3o�G6k3P���8#��f�t	ܴ��Q��.�@����/�J�;�S�>h�d�Ri�hJV7��Oh�=/Ԥ�1�kʂ0��D��U�ȴk�I.��,6���!���c0�oɀǲk�a�f|�1y(�+A\��K�Ы9�%�&Ԣ�H8dU�v?�3�~��o���b#F(1�0���hP&�5p�2���`/�ʳ�C�'T�����̰�l�A��۱=NB�"�v��.v��e���
ɰb�e8�<�����m	�m�C�d�� t�p��<%�����;��N?��׿��e$62�����3�f�.�8�!��;����Zal��e��r���xE�D����9�����$���1|ė={�����ʿ��0@\It�KVʅ��L6l�,�jA��T��	�1�`E�m�ZWo+�(`��#�ZU�(�*#�@����/�O�Se� k����A= �
B�0�wbڝ�{L�>�1��X�Cg����Q丵�/�Ӥ=H���i7|�Sdͩ����v�B������22[l�9TS4
|�q��)�/lU�*h�x@sV����W=0ddT�R�����k*g7;zNϡ�2�z���{�,)���dd�%ʽ[oאK�)�z�Itù��r��a�a�xH8f:8jخY����1g�UW��zVv�8"Q �.Þ_H��bdT��.��	CM� � 緼�M�w�K1��f`�ƍ��g�����4M.��{�,@*D�­1��< )	&���`b���1���]
ޭ�֧%S�@�q���5�46<�����Q�W���iz>���'b�`���@��D�!��@��Q n���xȀ��׽N�?�|M������w�yg�˂�Y>L>�l_G�(P��Ǝ�&~�	{w�'G[��I%Yg����r��bѩH���c#����#��`��}��zV��L`G�B�a��ˠ��/�\1*	�{�W0䫮z�zI ����؏!�XM�}�ٺ��k�y��3]Ѩ"a� �
j�B�rg$�Ŗ�����W���a&�)Kr��ae�o��W4�-"�1h0�0���m�f��@( �3�T���x���q,Ap|���~�#�aψ£��A6��j�v������M1�tH��}�谖zA� ��A��9 ~�J��\��j"����� "߬$R,��f�r�[����%W	Md ��{����1z��3�Q<A���J� �
 @�E�[F�# �XK��X���Z�� j�0#Ѓ j�'Ӌ�4�[�*�xܡ��ry��u�}����I�q�K��0U�/]>(��|��iш�1��64*��P�c{�xA�ш�1�ne���́m�5�|���Z��m�{��#���Tmd\JT'C��K_#KJ����J�����{�O?�9��iL�	�{G�KS�	M���e=����͐�-j�� h�#�[jcCK�s�Ӵ�fm>�I�'���'O�'*K0h؞zz���茡� ��ؙiob p� `#	��h̳�d��c�j,�+o�\R0��EѬ�x��	 CK�(A&qs7�x����4�%t/�@4
@I��x��2�)l6����l��m�+N���ַ�_��_u6�;�� �i����m<���MA�v�5]��W֟�/���R�nؿ����zc�lT���@��K./S�ll1jۙղ?"�#��ϕ��/5�-�Zݗ�%�dhDd�Hu����%Mx�[(��N�8�˞k@ژl�bF�Q��>�W��W�{���El!#F�3�[L� !�*$�O`â������r�2%������)���Z��n����Q�)4 �?�p�P5п��@���ҵ��I�[�:�K�3-S�Q���I�c��M�����5������w�*�x�2��WF��(��1;ʄ
��
"�\�B*�]�t9R�*pT<�R��0��g��R.��z�e��f�4��Be<	�e��Z��|�{���!���R�� G��2P��f5�[n�E-��#�T����nE"��(��W�?2d�A[S��xއD�Rr���& L�\�ׅՑمpcL���7�$P%@����K�.�m�&�=C������N�n�mG�	������n����\�����~�=I�;�&Œ+a�O?�t;izG���\���}�q��D����O��/ɑ��a���/�B)$KZ����a��1�RK���$�$\d��![�1o�!h� �Pi[X/��+j�t�������F���4@8����Փ��F��t�F��(�=�ܣ���p�`��t�t�̺q���g�Zb�b�v���
�\��������O�o�2y�������T^Օr���Q��� ���AF8�2�`¹�R��x��Ы:�P��ȑ1�η(O?�O�9o��
��QU�Y�J	p��G�3)����%I��	!���{�fDw�$�D�	�� -A�o&i��JX�]԰-s���m��(��t�����#L����F�����Ibv�#��IC'�r&�a�N�v @B�wG�@;����'& 3���3�����y[���;�1�Z=���4T���!����3��G���p��cN+�%�s���(��
�� %@HT߈Q�H��=���o�A�8��B�*w�X-�4��G�=�EŜ[�h����e&ۡ'�"@�`l7��x��A�q��-�o��D���t��'�5�ˊ��VR�l$	��P�	�	�V;C~z��4�����!�M'^����%S^��G�=�xiE�$e+�:Z�\���hM��ukd��^��	�F2+k�'4:��xE�"���\G��	-�M����)yAM���a)���c>{�OFd����_��F1��;�D��h�U�H�^I��m�I��u,��b�h<���`��,��[ u�+�x;���ΤF�i��m~�#�:,ms7�RLg���Sh=���Ͳ�6�O�lp���.�ț��Z9}�Js�5e�����ۼVPȓF��rѺt,����%cY�r���(w�����0���+H���t����a�Q�
ؖV�7������*�e���k8���m�4 ��m����i'������
Ϳy�������W_$�>_F���oH�kn�%%Y�AA]��¹��2]7K��g����Uv|�����V�%�Ε�����=�<%�m0+��`<�KO�Ig�
�)h�iE�:I�l�j�6���,�-��`ʻmwޅ`��9����Y���r�\w�I{���kd`�82:�G�{��F@Å�HZ��UU��Ē�ͽ$ryy�L�B��s�(��q�h.n��W�s��^s� w�X���a�}�[8����
3�b!d*�k�UO�U��pڗ�H@p�}@a���YҨ��&���hp4/tɮ���ޗ�S��}���+�'}��_;��b�X�#inkʼs���*���o�`�R���3$�>�TʮV$�`��nCnP��W�zz*j�����X,5UIƴ��I:n���$��L��|�$l��C���eɁ&U�hؤ/?���Q� ��G�J��%w��7f����J϶ *�\r9f��T��������/_�Ï"��z�R����.����H�>f��"�_xN0G�1\ՌN�Jq>e:㺵Js���)��Ubs�l!@��jvA>Ɔ#���5�����ȣ�J����+���74K�����D',	�p'�c8�8'¹��2�N؝��Xj���Q��P��[��CU9rpL#��9u�iV�������Q-�nV��Ɛ�m ��u[U���e��j'��Pf���L8.��G=��[�k�B��;�=�Tn.s]6W�G��U���=*cպ��`44ܐr�Wg�(4������)��șq./_It��JQr�a�%�u�ZS��4�;�P� v����n� �u;�-��خ��v�9[��h�ߵ��>w�I��LY�PD��$�,l$��+4��&J�-�I��pa���Q&L�l�윞�R��J����2:��˨��<�s2u��C��X�A����eI��3�_�¥c�Xv��oZ�dfq��S��d�K�z	Cfs.����
^B�ό���O�r14���{��J�Ud����s�շ��a�F�s&c�d)C�u�L�Ê��b�[&�aUb k�� ˀ.������z킟�1�EG�d��$���a��1{zz�Z}̀n =�.xhHZϭ�՜�ņFBR�(~G�
�Ff8�^D
��l��j�T;п��!8/R�m۶��}�X͆-� �cr�%�ȩ+��/c�vH
^Yv??,���#AL�k'�aU�\���[�	���<(x���m���_s����(�����JWπ����@���$w�nB����Gi����d���$��l Z�s3�Ta�c��8����-xEl���W���6�+�0�u��o1��3a���&��PNA�4\���(�(�2�#�rc�b�ID�����d(�<�c,�^���L��kց�I}���=��v�{v��Y�j�,]f�����e���X�W�è���!륯p���2�U\�9Qn�w͊�e��+e��k��2#��,�{�"8�l� �w<I�kV���s�	��I�ƒ��E6��DJ\֤c}8V� p�եy�H��w(���cH��c��"��� =/����$?�b'���E;˄����:�:�r����~
h�,�����9���N�c�[�7��;��s�g����Td3_;��L�3����s;>,6 ��m��dQ1�����|�;?�姊\y�y�Uꑣ���<ui�m�M������Aƽ%�s��\���
�7 ����i��C>b��3r�+6��ҵZ�hp`�2������Wj��昧j�Ł��^�n���oЂ�x������T�A�3���F�!���r�RG^x���e�&� �ׯ_/7n�ԙO<��w�}
�L��4���0���.��eH?WR����ޛ[z����Y�K�}E��,�UHB�Y�&���ej��$q2���d<N��$�q9�	�+�8,�)��n��lV�f�EK��u���Ϲ����{���,��=}�{��Y����w�+��x1�����ԧ>�0av:���ݽ�,(=̗]��{�2�=I�u�<��:9��9dÂ2�d�����`�u	|F��]�I������ҭ�}N�շ�b�W�SZ �����56PE-�k<L�n?ŭ����LZ<:H�ƽ����|��7��[���q3����t�g���n:vl13�L�23^�2��U�y[�l��:�x�С��]Ď
̴w����Jԃ	�b��|!��`1��Lވ=���ݟ��g�b�A���1�y��:��p�ȌwRQC�; ���W_�����%5��vJ�U/� Tt `L�|�/{���������Ed�2Z�������M8�ߙ�]q�tF�s�F��4�ޕn�w)���>�^�ꗦ=yw�͢�5҄�6ƻ^1F��~������=>6���o���{aW�0:rd9}�K��y4��}n:�A��Uu���@�Y�0�5��0w�za ���//�-�+l5�ھ��o-Y}-��|�W8R8C\��XU�n8U�w�W b�
��`Zވ��q��B�TuG��d�3���b�W\�b�B'���Zn�����+��F��1�bԀ#�]�a�9�
�dԏ�D��3ϝ�nF�#��i���Ӓ��V�6G����#���=�Kg��V���r5t�u�J��ԛۮ���%������u�f6"��jf��↶��F����%(������{~nO"���)������!zW�L)���^��������Zv�.Y�^ı�_�����fS�hZ]j�=צ
�R��O}j�'~_�3��ߜ&�\cm�
 .���.�����P`[r^ r��{��ǘ/�݉�s�}hV�P���k�413:">�q��Lci�%[�	O�y`�=x`!�����w�tɥ�(;�m?��T�^�P]5��_i���"��On���V���[�A:ppoY(`��$���bj�T�r����`�a,�{�����׿>�����9sPi~��/�(��z`p@�<N�9F�� �O�g �#<ª��ک�� �:a�Ӛ,hְ�o~�bE���������Y ZU�_��إxO)w/��ӹ7�x�D�s�e��7��嚟��g� V'lֵ뷊� ��j��28�<7;H��ޖ�>��~�^�'P?�:�i�5̬??�p!��$�ο͢S�-K.��1���[�Sth\��}����y4@F?m��ڧz��rQ���vjYԪԹ�"vI��F��4�8��L7-�׿���;��a������j���4�5J����Mb h�8�=I�UJ�ˆ��R�N�Yi��S�?%D���h3��*N~��wx_�)p��7��#��qb�y�0����T�h'l9 �w} :���x4�-�-�8�-��~����78DQ�?�y�+�Cf�!�}�����ɶ�K��H���_������M/y�3�����_�UE��'C�U#�;���m.ޗ^"�lKL��;n�N�h���X�Dd�n������T��g����\��Y?�T5~B��������矕�ߟ��|� EY�̆���I>p�#�-O�w���~����{�-	�N9C�DL?ap�ȹ�Pe�u T�j'�JǞ]�I |�q�� VQ��j�Ӣ��6[#
����J�{��Ep����=g � K�U��P������b{�7�]��r]�Q�����¹0���������ƸX�^�i*��p9��k^�Ͻ7ʹ3+~�<8{R#��=��H�J"�VI�<U���$b��[d��h=K44r���T�	&��]<z�ȸ������v�"������n�yN6Rg���؎��/��@3-.U���>Et�ra����*��!w�|�+�}�J	 }��^W�v�3k�H���Z*�b<� ��wU1�.�<&�%�h���[ �ƹ  �����������[�R���� ޣ> ���}���RA���*2�XE���y���<�$��KGsM ��y��P:��a7b `ٺ�hԏ/zD�VTX�,��XZ^z ���I���X������{�M�Z�8o ���/"ب(&��bM��m�yy.&o6'�);�`����[�IVϹ�eO�ux�=�N�� &��4���L����a/}�ۇ
�Y\^���@"�e�f�\�>V�N��M|u-Q���i<#����+��+��ha� 3��,�b�DW�6d�u�yX�ϫ�W4*y�5br0>7�x%�Vq���ye�~{�l��t�ܗ!|�H�´���d\��bu=�N����C��DM!0�.���v$�Gv籜���ă����u_��O�E:�A��]�b�L>W�@{�(r$��%Q� %jy��K�V��ʸ����E]�j�0T5�*��=M5����I����C��Oг�Qi��Y�}���p��jYXN]j�5g�����@��}��<�������ԧ��g��IOf���	�B��B� ��x	s� >��a����// Ѹ��_��_M��dòZ�$K�i���un�cP��u�߰^ū`��5��'-�@�a#:%G�ca����]E}���g�C���9�������i����.�@�f�
��`��ǃ�q�tǝG������ئR@+���#�	��E��䩨� ����ϝ%��z������"Fa�EdZ���u�ұa��i�}��Q��jUE�#n�ކ��M���`���@:� �Ġ����N_���Ro8�v��W���Z�J��5�m٩�8!�vQ?j8CB�s��$aF�I81V!��=���ʈ�bU�-%�9SU��t�[2a���1��;�t�X��JS��aEݬ��q���*������s?�sE����u����I7L��9 !�z���q�U�5h��ǎ.�ߙ�T(�D,/̏4d�͉��N5U'�!�
�'篛�����T9�хq� 6�kâ�@A����n��i���zl5W�ˣ�l:�o���}�53�f��i��+u{��U%s0 ���s}����%����__t�	� ^��/�B���K_��d=�*+s�|1߃8��*=u2�zL�w����T	�����fba~��0&x��߰LK ���/ܴ"1/:��A;Oe9a�Oy�Sʵ�h�r8\�{BC�=G����c�V���y9;w_a���ZNS��}[IeY�n35ơ��;�!a߸Kc������x={_3<�Z���?��	�vr!��>��p;�&s��0�ۿ�_��0��]��G{i���+���t�y&\������'�u-�p�*6a�Q?|�_,ċ(]���[��������19�	Ŕ4M,溚V�^���o�h͆���j��R�#3wX����������V�\X�5�!��%�_��&��:��"2��`��À�d�X75��XIaȷ�r�:�4�2p:�n�����b��G�s�:����k�]�9������/�M:t?.xc_�̊[�,�dq�2�<=����L�i����y��18�tD#��_c��Q� QU$kv����Ltth�5.zi�&��w��=�L��6S���XF�@���a�xhu���UWѥ��t���$}������w6��ką��&k"\7�֫�G����R[�w�1|ٙ��xo��g��y��c
� �|��a<�V~W��.~���RZ��I׿�����D������kj_:t�r���嵚�d!���R&;�ɜ0��}��������da�>D�џ����xЪ���b�c."	j�S"�?d̮9��\�:΃m��a��i��= �k�
h?��9�Fg�ܕO(:��sh����u��Iv��`���>|���$�G'� �)�n�p��x��_]������c_����{
�}֞�g�{ݖ��]�Ϧ�G�������q�S&:��V)-]�p|��8X�N& �7T��G����*0���,��~LT�i��B�A}����P�'i�L�{=>TU�QF�`��p�İ�hP@���gU/���	N����9�*MP�|���Q�V/��-���;�s��ϣ���B6E���e���ܳ)5����s�-H��<����@#�qv�H��;3Y�휛n�클w��|?���᠚�s��
��b_��hyȚ}e�-9�����8��:"��+[UltWaɟ����٫S�
��0r�1���c��K�诺�:b0(;(*�Fw5��3������Lam_��m���{'l��N+�M�/
 �VIgG�'�k��==' ��Qrq���:�I�Ȼ���=�%�N/}�uU&���|�_|�+�
�K�V�\���aqY��|���	�eE���=�š�Ɂ|�^���|�P�[6����~ٲ#:c�����S�]�)�9�ދL32Q�aLQ�u����q�J��#�T�yd�V_�Y�z�D�d?:�K.<w��7,A<J~e�5ת��kՃ�di� ��IdA?�d�3Οh�	� �5�'��1�W��x�H��習���;��u^c��kj!�3c��0����qǹޜ�(j4�o<�)
xUn.���д��է}�[[,%%�$��F����cc�N��a\H��^͋��΢��b�˼�E�/��n�_��0��.�@B�I�p.�n�ݜs�M硎` `����?��q�9�~��	 ��3�w��?������w|/���ki�����x�̍˸���p�*�{@�G�υ(D?�@�L��������6�}d�ѵOp��h��Ah�4Y�b~+7(��5Cb���	�Q�$0{?.n��D�n����5Q̶��'?���JUo�%���M�׍ȹ%<�����_�ӯ.��q������� nbq#s�� 7A��im�0[4r���Gy�U�����O}6����p��x�cӹ�<�����d����_�&m>_�SЇ��<�����@U'@�o�1@���ߙ�V���{^�_ԅ`��h�h�9U�bK��r��
��Ro�Q����93]����	(?���"�
]���O �u��7�u�v�s�5��l&9�'���an�=�9E���6l�Gü Wf�L�t�Э�ܜ^��Wd����n��(�bW-3qq���l4� �lP�0h2w�v�;��0�3گ�GH�=/}���t#�n8NP�;>cK�^9�qa�Ff�y��
�W��2�"G�vL;% �G��q�,�MH��8u�)����5"��ܜ<FՖ��(mE�瀯h0�*/��>c�37P����p^���OfU$l���Yn�;����,U�;��̀��S��?���L���� �H�3{��oHވ̀��Zq�g&ܠI"�wr6��C�;�L i.�p��Z�7S�!�W�}�1�Ҝ(�ɑFh4�K�Q���Ǆ�����ԙ�&ʰ�ȳ�FH�������9(�n4��X����R����\�1H�΄��Q���
 �~���0,7B��$N�i�w�f�4�.��QZY��zG��G�^���Q	Ψ�q%jn���ˮ����7�'�('��G?g�&��)�9�A
pH �}��|0�H�'Rt��.:���rl�L6&㤟�`6���`4�����S}�s�0>��0|��F7�� �|�����I�B��'HMH��ؐd�qSQ�%{�) C@���Z.���/�'j07�>ᚑ�sN�ec^k�+�����=��}�	r��n��e%�Fȋg�3���X���^��X��T��d���֓m�R�;@������R�mi~�=Q!��.�t����VW�\�j7��h�q#a���H+lB?#�b��ߌɾ�O$k )�1`��r3�|�K�.k�����i���=��	�pY��qb��Z$7��}�U?_��xy��ޛӏ��C'`���V^���O��ѿ��22u�V\U��.�-�.5���#�o��]�1?��47ߩvw\�y@�����]|K��Z�Zd�47��X#��%�3��cq�|8�`��=��b���5�y=@�	���sr=�'��1n&61�}��pO^܇@��`� ��K��T�6�,����*�(F��l�8�RB,�8��3D��碿8 ���>�*��d!r� Td��C�ٍ����FgF=;cʼ�xv��k�q�A�����Z��@|]��+7����^釾aL7�i����y���u�hlr|��V\c�H�ֵh�%�0������-_�tZ^9��W�TV�Ro��O%-�Š2�>��������L�N���$b�c�}�ܠ����\��܏���S棛�7��������4���Ä�P{ǖ]v,B��8=3��;@�A1؉�Z���� 8<��� L�2��������X��L�]�RGk�ĐBrZL�ѱt���k_���o?U<�٬�y�\|���xK����c��+�s��Y 0A<;;����d�y�(3��Ȩ��::`�o�0��bԡ�W'Ɏ�(e�dt�������E��Z�z ��4��� � '9�x�\�  	�`��Y����8��XO�7��H�ȸ7�ɴ� ��/�ʋq�1�[�+�2^�J�^\����Fk�Uf)���z�2q>4�,�v���M�f�,}�Z�J����l&|��������D���jc�(���u���^���7�Iǎ�*n��3.4Y�_cCl��h�`�C�����9��l|�w���*PؠKQ�<2n�ĺ��2/�|�Ӏ���uPI4OGe|�h\�����a��Cgk}&�{x ��i@Y���q~ݓ\�.VZd/��5�e�F �<��n�X�巼8]x������4���.�;+7"sX��D#���a��g�0� ��A �=@�Ŀyo Qt�t�@�
:��d<����u�q�0q����@�_���7@������)++��α�ȸ��m��c��
��: 'ǨnBtw�	�	�@̧Ap]�	аy���>�=�T��{�ч,n���o,Z��A
r�`�m�9�
�G�c��&2�ڜ�{��$����w6#E�`4P�M��J-�M���dW��#1���m��7��1F7S	W��O�Of��
4�:�t��OM���_������ݗ�^N�),���3�ɿM�յD8�$9Gy�����$��x�zt���s�����%��8�W�	c�ԤD�9"f�~��eW9�v���'��ڤ1�&�L��Jv��]}��.R��04���N� �N�\����H��ufK3��dYJGg �<#�kp0�1u�<��[�d��hX1����So̱.>����j� ñ���KF��FR-� � E�n:>���cf�WU-<L1\�~���Y ���L AF
�D77�Q��T8��D��F]8��Y@�X� �̒��&�Qm{���g�"�2H��	�P��Fù ^���D#z谈�
��G>�w>3/�~���s��K編 G�����������@�7� :�W��Fǎg	e����=��I��{Rz�eOI��q8�%(� ���u3��z�5{�@jڏ<���{�n*V��Q�F��-~�M�괂���r�Y_E�����;���71Z���X��7ͤ�c�<yVґ{o/,xi�P�`wםKiϮ����V��-�T|�["�.�BTsL��04&��� ��,� Xu���H��Tt�R'U^[�'���ٟq�k��ا �WG���ʱ��\�c`|����s��Z�Z�#(��k��Gi�DyY$ �U34[=�Ϡ�@����ʽ�QﮇC]�eC%�􍢪9@3�2 $�����k���`7�=)��F�8+��-�:D7P6DI���0�w��\^s3�3qٗ�{9}�����9���RI����!=���46SoP�0X�������h�٪m���X����<Y�:U���	��E��J���^w�W���xF7��4�I􈀙�K���.>�.��|��t�m��UG�u��ؗ~x0FB5*�Y�k�=K]Ɩ����+�5	\,,,�	���{f� \FE7����䥩/s#�ݱ��q�����
U�?�������q������ת\x&�	��S]��e�����P�%����iaG��Ёj(� #�� r#]Ԝ���mi����2���ߨO���@�uݬ K%#��|����W\1�ce�@�õ5������_�}���;679U{���k�ԯ3sԞ��J?����P�;�+���l6ͥ��=�Oyj:�����-�O�Ae������Q�3��~��\��8Y�\��hC�<R���g#p>m�9��6��Uҝֺ]*�������؅, ;�X��3Gv��r�{���ߕ��⢴�'k���8�5>n̂U��kTV��+�0W�A+J+*��M[ɱ,,U�|����vk���;�"��C���T�D��!@ �y�� 2T��H�� J�h��J0�����Q�j?*N�o��c`��b� �1�9�}��9@��M��{�e�</��Xm����,un���x��Ϸ�0��o�v�zэ���=R��� ��g>c��yO�rO܃���+����mie�xu3��ՙKwޅ��0�u�iiq%s�,��D��_M_��;���O��*�Oou9u�k�ݴUD����<��u+6IQ}�D�9n�_�P����V�Ś_��q*t�悎�Q[�f��j�	�R�ޏ��Z9���n�ñ��ư��2���x���ΕdR2��;�LD����H���}I��E	u��'lN ���Ɇ]��O5@�0Ѓ{U���q�����p��waEi)�J�� ��|n�7i�.�2{p֪���N���e���Pk �|&+���>��g}J�����oA�<ԧs�z�"�s���_�{g1���G~ �㬑Q��:�is�TZYi�@�k2��H��k�lg>=p�p�x�ymeIs�f����q뭩H�7S�P��dY��{^/�;&1�cں;�6<�>�j���CٱQ�w�����hQt�܈��)z��]���w�?�>��v���ۊM���͋t�'}����ˮT��UڞQ�r��\@,���F��K�]��_�{ݗ�C������{�u��g��M��GР}m#�	���c�e�@�H��]XV� �Ȟ�q�Y�C�X]4��n�V���F���7���]m6*���ٜ 4@��ͣ
�ee��*[�?���+vC�9�q�T��=��<�c�}Y�����97� �q����g��8�\�f��'�u��%B�7���AZ�k璟ɛ,��a�V&��iqeX<%�>;o��"�s
��5Ɖ��/nt�s�"^�}�@=��u����I�N��Vmk�Q�7�r6��Q_Y7Z�p�e�N��q���Rv\�?J�P��ꫯH�w5��0ͤo�ݽ����+--c��)���l1QRe�{���X,�7%I&&��hp�K�j�c�O �jl
?�:���M�P�F+�6Lӭ�H"��d�|�ƌV�D�@8q,L̠��	ȹ��Y�d���� 2���Or��{�J�O�HI��
2Ґ��q�:�ܜCC����;�99��bf�������a����>�zƠ�յN��^.1/�sϡ��q/2f����y��o����d2��F�w͑�}%�⫟�^�����\� ����F8+�uj��ހM4K���q�8#Q�g��W���؅A��&���}��(���	��)u� <�'Yv�F{,���+���޴U֣�L�"���Ț�nRu?��8��1�W]�_WV�r4O�t�y{Sp$�u���{:s�U�fv��"Q����Y�k��i��gq#�i��j
<7� zpO�v}!c�W�u��b�w@s��Ⓟ�j&Q�xt��h����LQ>NJ~g�f܀��70<�w��ƨ�t��i�y(�4�Ѧ��c���{NXolO�1X$����iج�5��|��i�IT�9��3�a�ul�;��^ �^ݸ.���q�D��g��v �����!Qo���XIg�1����J����=���'�o#ϫQZ<�(�`��crS��~�n�]�~oJy��<�u��@c�*?U��,�����.�{��%Ap�E}��w�G3�^�1 �{����w;��0���F���#��ZlG���zb�]`u�v���2>]��M�ڠ����{��(�w�Bz��.K�����Ky?�J�'��+k F���*߽U
Q@@0S��ϲ�Q<e�I-�ɈQ�b�f�p���Km����n@5`�-�u"�J}��o�i�z�&���N�E°�wu�����7cqu2�9N��bۮ�9��4:�ˢ�k}�5��G�l�C�ޓ��M�����Q�yZ��G��j*��T���&��������:P�p�W�e��m�=��m'&x���.^Y��6�����:��e n5�A�hI=�və��	�Չg&"y�v��w�F~;�,��h�(6hx�^W?΍�]Ռ�O�G�VW�Lo��^�~��^��ҽk�;R��0��󰪶<����/���K.�l4�ϚU�{dN���k����0����������2�4���߭�[\ [o���������A���e�ݴ�nv���u�'�L��5�	�H���l��¥�L#��|�ӟO��ޑ��I���/K�?[ x~>��X&@�����	�/�wd���h<��� �$��c����mc�e/��ؤ�9�!"��6a�m�j��G��(�ɮG���&vH��d���F����n����=��\tx2>E�1�ц�H��L��ٕ�{)}�c�~��ǧ'�����xHL���y. b���,�Z*�4����]��x��x�C쿸����"����xYr<W��~Rډ��F`u� 6��nv���Zu�����F`_�~��6z��4��U�l���0?��>����wI��L�=�?;�R�#HPe%]7Қ7Ud���X���J�UPۊFN�EI3�����|����͙m��{)�C;:�̄��l��`[c ��y��C?5�;{�7 �X�aS�?�u�և�
02߭�u=My�0a/�N���O1�x�:`AM��s�Y��W�����7�M�K�4�!�CO?Uي�ͱKZ0Ѝ6WG��U��F�G���
S毕�}���$�ƈ��KM}q���!=���=��6E��g������`i[�ش{8Q�?۩0�킿�4ͮm#��4��ζaq�Dm7$��Q��������3/�n�B'Kγ��[J=Ԙ���iϢ���\�+�*��Y�u�F��f�+mp����_�fTc��*��k�������;�AC�`X�,�kT)�V�Ki�W�^v٣J�E:�/���N�E��� UQ�&G1�.j�26_�-:����Ź0��c��q�������/3%z����G������´ɜ?����Y�ze�h�Imb�
�e�5XV�R��s�S�z��'��rpC�Z����^@W���&�h��3��a\��Qo�O�O�}n����|�����j����`l#��Fg;s�e�o�JDe��(DXE��BԯJ���8�1C�����׾�����>������+��h�ǥi��P�{R�^y啅0�1u�\��� 1 O�KL�Ͷ�)��v�QF�E��2��	a#�ݳ7=�Q�MO�3&��`������N��YB�2�X�Ɇ�\w׏�����p�&U6�bt E�?��?.�jb��Xbm��ĿF�'$�����^���s�={h�~�2̥����ƨh�[�[���L9W���`�L��4�Q|�( ��	}<�~�
���a�s�2���I�Eo�6���7hlv���Է��&��9��t�����O���uY**J2�eN���ۓ^�/H_���gr��slD�Ƽ�g;%0jee)���KC�;���\M!��iQ�F<��,�ɍsL�)��X$h� `�qx�@H��v}qM�#�]?�9�)XCRx�m�JH�`?�ߝa�@�/���xEz�S���@y���9���� X-���z�K^���O�tRa"zV��Dڋ����u�1���Ό���>s��6�K_��t�����yr,��ե�UP�F�P��p\�5�b��DSfu�F����/����
���e�B�-�4�<�����RLS�._�z����'Y'|*m+�jlu={�|#�矦���s3�]7����a�Zy�o�
O)~���	 �ٵ��qՕ�w~���S��t�E�j�H���
��t�+(e�x�i�z^�a��3�� � f�j�pǊ�G`��W_]��
�`m��|J����{)X��1�馛
��}�Cw�v<bn4LFX�O�9�I���?���%q�s#hS`f{� D ��l=���� =P9�ܮ����{�yt ��}(}���ۍ���"U\�z[o�\�B+U���׾"���t����y�V˥�܈���A���H��	Z�6
;��U-T��GU�F#�9$��琨_/�b&�k`�zf8���g|��i-�F��'�m�з���TJh�����ot��x7A�I����rNKKi����[�>��\� �c��ֆ�N&����Go־m�b�#�Sy��J�:�=�;_gO:Vr��t��/J^zA����b�[]=���K3}���� $����Ӌ_��w�[5@H{�;�1I�dȼM&R3�������;L�B���"zd���/6�I����a¨#���w�V������Q��С��y9D=�D���H90����t�;m I����e/+�!₺S���O˥���;jW:���F���oݖ�;wEs9�J��]�����g�9i���q��x��/c��z��������\��j��J`�d�%�ƅVw@����~ְQ��,t��ͲNG;ϣD�{��xZT��bܘ�<Z������77b�"@G�����M����F�q�|��p7������~��<W���=i���]EW<U��� mU������ �?��?+��@L�Ԙ�Ԡ$��T �%8
�dyf ؠ���գ��z��������Q�vm��M��N�Ǔd�ߪr��t����
Ӣ�0�J���������≘��c�w$���~��������=�yew2��:��ӛ�[Â��i3��a7����O~$?ǝ%yLw8 Bno:t7eY�dqk0f�c�`������B/��Xj��b���gdr�䜗�nu�1Z��_f ����l+]������~�3ݝ�h�L��T<�@�b���h���+螥Ǐ�o:��^O�Y�:k�N�
M+�d ޕ�����#�#7|*�������ƹ��O�:�y�i8GC��6�A�^%g�)"�+�>��t�7��X<;����s^I� /�����D�Dc��zt����<��#���O~r���k�{O�O:�7;��Ǐ-�7LG`y��7h�.ߣ��0�$�7�	�����s��a� UX3����ԸP�b��Dy@x�A׻2�=^,��A��[�,�lwW2J�;��z�H}���Dp��P`����cSP����CYYd\����v�m3C�N<{=�JF�/:���M4_O:�]��Cg�9�c��=��!�y����������yMt2���Ez�kϧ#�g"p��^�x����Sk�R����Өt��3aUeJܣ{Я�گ��O�_�ksx󖷼� ����rN}�G�R���g�:��F���H�@`�C�Q�BBQÊ5����L8��Q<�IfЏ8�s���&�Ao�>���6���` ��P(>��3���ท���e��X:�����{�{Kgt�����N���
�u�U&%9�3C�Q�O�!��!ї�ۣ[3�g�|Ƥ=��~q��|�I�j\b����g����1��� ���!?
��V����P��7^s'�7b�H���S������77�9,Xi�;+�u�Y��$N�y]G���:uuDQ���Y:�f�^�ղ4��n����i���k���-@�_���&x�j'�cLpϽ��o,j�c��g?��x~>ӥR�˹�_�
�f�i���4�D۔BL���&�W��6�U`o��`�F�?Z�,�,����������l�UԈ�~3���b����`h��\Oy�Sҫ^��I'�[���N��z���]��a�:"N���]>�Z��,n�K/���ӘOݕ=yw�?�g��#�
�� <J�zz��|��؜@$]��ͤ#�� �A�z�gN����t��$�}:��MR	.����3]'Y3,~2���5ZCD��l�w�D��Ѩ|�����M�fb�����Yo�Uo+uB�Ľu����8s�T��hB��L������g_���\,7�T��1�s� \E��<��5�����t�5�U ����T��?Xm�g׌^��4�=&��:JVR�n|f�cQ\pW��Q�qj	�OHQn�^1�IRv�V��Wr�iD���b�[��s�P�3hQ�Q �'bɯ�ꯦ����(:|����g�z���4�M��bzы�Lg�����-�fs>�����?�'�:��j��W���/� �Q�$�9�>���V#�d'Ϧ��	�,�v\h�?��Û�u�T�
�N��9��֯����1���T�*Rm��Ҁ C�a����H�G������P��������4��/`��be�8���h�jN��ʀ`����tn^Co���^��g��YI�n�v�����l����h��Kq��\�'�nhu�6���/#���3D�����e���7}�zrܢ�>������Q���4�
�muO�7�n�5���kV7�5��wח{l5��x�~Y�zN�ĺsˢ-?��w���\LX6L�-�V��!�b[£R%�9���ܩ��E�Jn�NZZλgcWIFR"{FvY;m���m����lOQQߡ��1�}�p�~����QT���
F�i���ТԶ]��@�o:����o@�o��
�3E�����ck &��1��s��� l�k���y�?�Ò
��ꗴ���R^G)�;�.�i��N^_�y"W�(�����̩0�q�Z��(<Pi�ˢ+�U]1�`8��e�GOu��F�K����@�3:H�� {su��5[�Q���7^̣�I�JG�@FQY@�n$��Id�E�b8���Aa��/�忤�����x���S�{&y�@�p�}?梒�w��]��G�N����R��Z,�s�3%�)Y�ƽQ�xF̬yKl�Ec@l��R��4&N�i��?��(��F ���F��,+&������i�#��?kL[7)�)���[�g�f-���5%	2$��9��"o�����N�� ;�y]3���X�Ъ�Gp�B4�q[��sh��(#&��
 f�*"r�~i43�����8�7�?��R1p3�G�/�/��/n�b���/K�ܝJ5���KH�s���&8a��qݲ����o-�qG�x/j�4��{��__6�?��?�����T��E�UF����Q�i~��I
c����j;�;ɶ�N��7��(�����e��1��y[/*���w��99�w�R6|f�Z	�X�%��������b7gpaLl|S p;_fASE�:f�i��n��_�n�t����%O&&��4d�..h�qhGs��;�����@�Im��;����X0GНi0�`L޽��آH����4 ���z���UND'�[V7o�7~�� s���Q���4bT�_nhQ�S/���@$g=p�qtKs���G�ܕj��J$�)�����.[\<�n��O���7~/����ї]����/���5���R�s��� �e�;�=�)��ozӛ���jbw�"}�Ā4ab*�[G�n-� �Smj$�����)u���	�����/Y�mt����,���=�:���ݭ���CE�a8L���U��������d춵�����L���|�L����7_K��c�׿4�y�A:T�s�@����}I<2S�Χ��f�+Y�e�yY�GЍ%�l���nH��F]�|i,D3ũ��1(�D[�}Ǘ�C_ɜ��1Y
I7Js@ˤ�}�g� ��Cp�XT�1�Y�}1�Y�OՄ*9ƈ�8/�G?�u׵���GԵI�3���CZ�d"���f5}�7�C���y��M�3Ӡ�7�h&1�RH����Z��d������Dʰ"9}������whх�y	Vq<R�D�9+fG��͚��`�5�8�n���΃0MŽ�ą���yl��{�7?H5QxX�G��N.2` �cd,�6>�*���]�c���g��GL$�	��\�>TvI]�bL��ހR~7K���G��_ �LY��~j���=UG�\�1~h�QO�99�������E ��u׶�g����bFOU�=����dT�O�G�����kxV}���KSt�~������y�K�[�$bb�� �R�����ѕ������
*B4���'Ԋg�Lj6f��Z���������轻:�\�2��ۈ����^��i�Ա�y�$ B����}��.}�Z�_�7X1�d�a���9�:s3f���/Y���4c^���q����Ou[;��F�q
���L���z��x�v����M�f��e�WUh�-�����>P���y!�DL�/|�El��8���7��t�'?����L X1zb<30�=:\g��:��,���`�i���iq)�`��=�@z�c&�gH�s�ʢ�f�Ԩ^��S��2���/�7�c
O�l1'(!��[��\� @K�����o3��6ꍚ��µ`�0.�1� �p�_4�>M���`��nP��Ju�lWM�l�����cY�(�l��Ak@��Nj7��L;R��	/��#.97}盇��b8"'L��Ȼ��>�id���ɧ\�Vz��_����� ,� ��9zaT�GT���i�/ǰ�+��`!T��4�G��	hƏ1��p!؅���0��lХ|��0��۱�^�w��~���(a�;��$#�����N!β禠��1�����fq��Pο��o.�9���hX7���-�F�6;�L�\z0��%�N]�_� ��f�z���{q*蘆zrv������C�YZ�1a�VRIo]�L�aEU�V�a"�D}��1M*c���<��s�n����-O��'���p\�HP��{�~ ^��^�xCf`�J��LMu�L�>�m��舭��� ��֔���r"�=��g=�n)Rz��l+�3��O/~�u��dl�I�|�h�
o��TI�k�Kq�:F��G��!�}��^{m��AU�O}j�p]]:}��Ma$�%�C�s^/��'�8@��%�N.���oi��#(�93����ц<��?���{�t�ŗ,�?�V�Šk8q"3	���X;����Iq�1�,nM6��mq�G>�ѓΨ&{�zhL�ed�X�|����W����ͦ��}LZ\>�fڳi�t�T%ܝ<�*#\�3��2�*6�g�[�%��1b�A
&2��&d�ɞNT'�zz<������T"����d��O�C ��������@4VG/S G�!�Vw�aql6�}�dqN��kV��5�� vӆ�T�ek��Z���'y��3�`�V��g\�Ĵ�ey}��3�<���#ŧ�����������I}���-0��V�@y���EE2��&�s���֞����#5���������;�#�ӯ~�u�6�p�����Ύ��^&�jeG����z��/|I�ǗIȎc�"��.8DU����ތ���G>RحF#�TY���/:����4YX��D���v�)-�.����%鬳�(�t[���N+˽<A��Օ�0����үQ��l?���80F2��W�i��f-�" �;��/-���)���ۉ�~�w ��5�(��<�����/��,Y/�!kG]vd�����l ��p�
�	�d�l��j<g-r �=�����:hʹR�C����l/��XI{����v��鑏if�r55;Y:Y��n���k��j��ꪸi�o#j�L����!pT��y��5���y�hxv�XHϸ�2.�	}��a�V�Q�~F�ÆŹq��5�Z�C#�X=��L�֘DUU~�3c�gb�`w�ywȆ���*�� �b#���_�bQn�� ���7t3�~���L8���Q�Ϣ6魎E�n-�����ay.e��a��׿����oڃ<1��مt��y@gw�!���n���+nzD�u�U���PoV���{��aA0A�ie�Q|*�������7��9�\�C"�N7�	�>��O;���w��2F���	b/�k�˭���K��3�p`�Jr���Ƴ���1�[/^f��.9�˔�fb��X��E������' X&AA�eʅ�f�`6[���0K����3�%U�#�����|��Ԟٗ��=P�� -�ߝV{˕zb�Ve<��^!46|�� I�6!0�������4�K�����
!Τ�%�i)CCntd\�_^0p���w�l�������k���qI�CU��7*��X����0꾜:��a�kW�zе���"��q����%ȸ���E����X7���a$ ��濺1���Ci~���*��O���Jlj�˱�i��Rߣ�����Eo@Ft=�FٝhηXbD㿑��N]�y"��^Ի�7���=�O�`gp���@���FBc-���%`	%����u��ArU�l�w�u�T��F:�z;�t�x���D��{����Ꙇ�� �p0�ڙ�\���ff| ��MeW� �������6`�N��7���FĜ���&��aM:��T�5�$�[p ��CUi��O��ԙ��E��������9O8d�\�v!>�3���[&��&�| Ev�<t��%�D��u���ۛ�PT�3 �;��z��q��p4�}�����O��9��Q��=�A9��ü�������
�x�\ԑ]2	g���Dܮ��j$���cܙsQ�|:Z]']7ј�z�0�!"V��l��74�&4#�8�u�� ����%��M窚EI����>��-�G�>��^cl:Yg��]ψ��TUmW{���3��Ŵrt��9X���_��-��/s�V�L$'$���� ����-�;�o6s@���(�<1(E�� �IA)Ƅ<��qyŠ��n�Q�9��G'L�j⍳菂�����swpM�nn��6�T����h�h�����u:��	�P��j\D��������i%���l��#�9��V�$q�lU��A�\1�������4`����i1
�D|��jaEN�4�o4���K��<�Ws1_�����orQ}�C�S�+�3ݫT���<��=�C��=!y��6##�p5�O����I&4�yu���J��ʌuZy]f������R�]��vJ�!g����J#��-���'�U��>T�#TI��FP�n�5͋F_�hߊs=[O�m�;���h��n��\��ϢU���-.$���4�n�.78�fLL;�D��5T�pK�/��u��,B��H���^�5O�cu�-�5n���n�R�c)���?=�nէ���P���;�
�űӛ�;�ft���m��H4�,Vw2��vԅ��Z�Z���)��1��(�,��*{N^��#���6d���F��:��sˈ���gh�����k�K�]rNڳ{��Cbڝ=xg�Ӯ�*�{�y�T�k��g.�������ّ��b���t;�y%�?ٱ��J�FqN���ʃ��{�T6���|�M1MuSh��	��`T�6֘Ҵ���\����J,�W�u}�h��u���&������G���E=\��h)=��'��g��r�;��sF��H���?�n�-R@��xs��19�9#d�Nds}hMvb���vYpl^C� ��wJ�q"��!���4ؔ4~q_|f�\��F�ׄ��t�ENc� . -���2Gn[ �ngQ]ǵP��ր	��@aY�(��&6��uy%��e���=���k�s�{u�(ޞٓV��t<3�]{2;���\���SXtņGE_K~�z0�FW�W��r�(J]p���TM���)��,�.�Ӣ�'��t�@����Iw�N�G}��wu�R���Y@]����ˤ�R���kO���0H� &���Iˋ���=,�<)�ͦ��F:|��#��w��f���VTaT��R�A���ޢ+�(7MdU��i��3T4�L;��]���玢*M 0o�^9,t�$��F��u�ܵx'`��ݤ?S�ZA�y��#�ٺ!a��/�fߨ������G�5�]��/�^�)kp�Vj��_����)�0����J:��FqUC3�j�O�+�t������L�=���cX���5�)��Q�ZR�8���������M�c��c%xu�1�6�Y���{-7��MAx��M��z�3�)n_щ^qJ�(]�Q�'{|/��3���Ȥ�P;�	��J�k�K��>��򦏦K/۟���G���۝Ť����®�<��lK������i�I�PWO�uc���i��Ӫ	�Of(�>O�q�~u���z2p|�ȯޅp����`�F��o����� �!�%�3_>l�	U!���u��X�����6"�h��k����:Y*kfiq)}��_I����ӓ���t��Jǎf��ٕ�-��(����-^��Z}�~ҝ/�O�F�C�_�?�Ҳ�$V�u7ʺ5F;�T����n�:����RS��-��Y�hQ�R���5�s�~~~�e�^;2��ǧ���Z�TϏ�i������t���7қ���~�.�g�yR�������Faヰ	�~$���|V7C�� ��d4ҝ����`@k��D���TtC�'{O�5"��m�2��$ǉ���A��n"��`%�B\;4Y6�|��*�~�<�$̣!��;TlH0������'kl2y�`�:��bجW���g��+�7������}��ON睷7u��|;����'�Z�*׮䫞s$�����9�;��ű��N�w���:j�5rwJ�~S���(ߘ\b|�k�_q�h���q�(Fx�'��,������_��1�zu�s)�=�O�<I�����&=�W��>��%���2�Gg|���Q��x4���N8Z��i��t�<W��  f���������<��w���Qw͹�zy-�g�C��Z�ܒD���Moð���)F� �sN��P�{�X�ي��:eذ�]"Q����Xj�Y9���Ψ$jG�<r�h���8�Z��v/��V�3ж��LN�G��z)j'��>C�=U<��umu�`���D����'8�q<tџ4�Tf|0;!VM��1�Zd�3{��^p��:u��|b�M�RUy��,�u[閿�3-/Qv&�R�S�=Wr#�$��I��Q��Pn����H����.q'T�m;�[�,شE��N�s�r�df7u��j9ݩ`�օ�� f���� ��c����9A��djzr�⼀7��]Y-/Z]=8MT��o�RN=zdt2;˼��b��Iw�u_&7�t�E�|+�ػoWQS�
��-k��N�7Zw�mbE�k�q�k�uf<V7��)��MA��sv�dQ�ڼM��`"�	±	�u����ؚ�q�E����w�-�r����R��f暙)�"��ԙ���"���3,Lx<l�ᜰ��u?tq4�E��rӌ��p;-2���9��4�Lk�C-�պ�wBg��׼�ll]r�����a���	C����bXSg�a�k�� �a�a�oX��Du��wDɡ�`�@%�kZ�����Un�Ʒ�$ٮ�g��m G@���5O��y-�:?(�H�Cz�fk��+�̠1>�f4u��ApZ��>#�����ql$�Q]�mLQ��e4K���l�gQ��-�.*�xg����c���n}���3�����T�k��,#���3��52��}/�ڛ!x���K�����t���ґ��y�P�1�q�[o���w{�b��v� W�nd�Vգ�h\U]��X�!l�EU�j2ϭ�D\n(�\#�ȑ`a[+`����9 W�lh.�h����P{L�8+��p�>�&��I�F?�Ra�|+��g�s�>�wϥ�_��t�p73�R�����JZ��`<[�ёw�0��cp��r3 ���g7��X#1���љQ��wx*lxsn������	�t�2Y�����|ŉT_Q\����Z�U�#G����]�RG��ܮaz�k_�.�p&]��+������r�s#ZM�/�r�4O�S,)��������� �e�i5Ĵ{��	6�	ڨqO���QԮ���4���zO�> K�Q}Q�����OY����wo�(Po�$K�?�b �k�G���f���Ͽ�{_I�����������lvP���ٚ�l�\��4���>����>'}�w����URY���-��J.��z����]�˳ҷ�	�9��a�
�p=.^�q���MAx8h�0��0�:�x1)�Ư��x���6M�+�C�k���D.ӌtu ���E�;�^��̦��ܚ�7�^8�Ծ�$*q2ڗ�7TK�>��|�l������C��h]7L�	]d�&Y����4釶���ʄy�f���}�<��l�uт.�#ޏs��PQIX)C�<���Vu�=�#�9�I/%}���h�,}1�2&6[5���n����O��s��tB>_|zgJƲ�\�����ݕ����Һ���:�J��]y�<��oN���E���$��.}�O2��\�`x�x��޴K�an&�(�`7�N��5"EG��O���/�[��t�f�0���AT"��٠l����h^O|��5�\S�g�'�(͝�&��*<͐T����~�+_O���L�+���);�K�~����6*�\)�R�yTÛ�M&,�g��o������IFK���͌s�xND�y"M/1�Ĭ��ɫb"��PĔ�Y������`�(���d7&׻�K�{%F��K�ϴ�i3���6�^&+�O��̂WZyø'}�K�ʠ|����p.�ʹ�{��t��invO��-���8^��h;����������I�Y���s2���<�a�)�S��-t�Pr�.+!���j�<��^z��W��{Τ�9�2LE+�3������:M7�tS9>:��>c�����/y�����t�UW����-��9d����o/;M�B��}|�����A���[I����Z��Z,9���y"��Nǎ؄��@�DZ�Vs.�0e��P���x�p�er4� A��^�<�����9����Lr��i3�>��O;6��Ģ�3�+ L_@4��i�\� g�,��E�K��G03�}��v��Jȵ�t����B��R�'
Õ��c�(j�Z	�ڿ!`��"ޗ�8�_��{���tÇ>��A��I�wq��OJ��|)������)��:I�d���70���^���� %%�ԛ;M�M	��4�~��+��#8w�7g k0��G�Z�CI$��<-�Q{�h5[�����)�1��,�'�ܓӳ�y]ڳg_��ٱa�N&��x �EN:�T��V�K��V]�j��ԔBd�?���.ߛX<V��X�1od���|�]��d�{h�Ҿ����f�f`����nx46$4�9XmuD�iup3�D�&��n'\��O�\UCXN����t�M�T�V@��  ,N6ve��*ki{uۀ  ���+nz�����Zt�����PE=�6K�����Ozz0��O�ռn��u�Z�MGC��s��u[fó��S�Y�UW�K�Kl-�{�/fD�oc�SQ9V��&�8S\�����7JV�x�3������k�9&����=8l�l����+�O5 ƚ��5��d�A�6>���yIf�ץ����j�h;1L@����`�щTL%3�ᛑ-��#�9���`>N\��h� �3�peۃt�H��bR^L��2��8��9�x$�#L�1�-7�J�<`�n����n�r�	
�7bB%��E)�%�j�ZQL��+{�0����^��Έ�6a���(�\�����8ǔ���0������?��-",�Ρ8m��lR�W=��'���[�HEs��H�����3N��B'��%��WRZ.��о�v�=#8X�a/-����[�y���+éj'��-�K���������x�;J?�[���CC�M�o�q�4jL@L"�9�U�P�tp~3F`�VQ8�͕�v��d���i �����~#?��t�W���~=���3�;Zyo��I�P��s��-�Z!��>�/y�K�w��Ǽ�u�+���b'�X��0�z�	�$�LN�����GfJ�~��-<����S+l���TJ�4LH
>�A8�t���I�	u�y�K�9D{栬PF㦿�0M�\��y^�E����cX��0�EC4��ҏ��wu�y�GI��晽v�H�k�Ɏ$��௚�r_���V�r$]x����F�T����.ܥ��<&u����/�{������ )�fc�!K;}�ӟ.����P3��1�>�&��� 5�;*��1:ڊ"��g�������1c���}n2��N���h0��/�,t�W����)`�t*`�e��{'+��Э��2QM�����:)asF�=�O}�:Jv�v�Xz��H���I���4�����ݝ���/�Gjj�	��!J�V���|����{؉T3>��殺���et��Ǩ�nX�fF���h�Z 0aĬ�]�ۚW���7K�RSVE7W��Ut�C��)1'�a��sG76��Dl��Z	�5�܉��s��RF�f�iv�\z�/�<����N��^1|�;s��qX�\j7����uG+�_���n�ES�B5�A�1}�я~��R� ��RmK�q��� ��
��>�s�^�(fx���3
 �G�h���X%qzK����R��L������!|��a1 vI� 8�BG;���� ��yk��s�k�oD������_ˠ����[�^L�������<@�i+���{�&��K���RvTJ��Gm ����H �0�y� �9����3�h,66]Æc����s�噙��!��t�YG�M��:\�M~���]�Q"�𞱁]z,��F!H�w��r�2��N����]��^<v��/9��~B�������L:v,K2�nI�ngf��R��y��ݔ&�rm��7 Q�#ρ�FX�)��4�0�h3�����
=�/��➼4�2���ê�X��;τ�VAv��^p�y�#��~XtK�nR<�)�5�#D�B=1��,s>����ꜛE�e���zX)_��W���J�]�1@#����X1��=������\zFz�k^�f��<p�8_��I�L�s��@nϰ���EO��&[cc>���U%�x3���0K�u?�m���h�tB�l��>�����@+; s�z��u#d�3���"F®)��ҪM�T��y�7��Bj5��K��0�/9��I��,5馛>�>�gQ��ЏN�3����?���l�uE!b��}G��׿��E%A?��.�U</�y�w��]�>%%<�x�3 �/�P�Mi���Ҷ��8��q�]C(��
Z��q�y�s�����bqgh��}��W�� ��Ibuc��T��xH�-����B���qC{�k_[vA���t��t�;���"��qq���2�.��#�/��>������;����oo-�r���L�1�e���"��DܿO��Qׇ���ԍ�X��X����I�J�,�t=&;�`�Sl�ޢ��{B�C2�'��em1��x����~�1�&M���;�K�X�a��fܞ��z��L��+����=���_~�3����ҡ�{�7��t��{K��fs6���R�3>-����y0ȿ�e/+��.��oxCynt�|nE��!�XHb�b1(��(�sn�EyN�Gm�=�G������ڈ���UG4Z�ҵ�[%x����$���ۀ�$oc-��;��+�1������"�y�~����������芟��g��e�q������¤�sh����ӝ?�7}�O�:��U�K�>��H�b�+j�F����Uʲ�Fy�7i�Ֆ�"��XMs�[��m*)���&���b�N���&�Ci�~ΓY�^G�k�s�qm� '�I£
�{9���K��;2��
�3�%�Xa���`�,q}��XŢ=Eo	����õ$@T�"�a�;��owf�sdm��U�������t�������aw�u�T�f��3c�W�,�	(�̪��G�e��������˛���"��;�,+��������x	YS��O�~�����S��k�2H4�L���8����'=��PG�G�V���ʺ]6]���k�ݍ��S��dwٲ�_d
ՀV:a:#�C��ab���\^ӿ�ɕ돆ie9�C?�/��<IF��[�H�_p^>���� =��\�u�-���+�? � �Rg�?���.̦?�fA�U��L��۽׺��k1_�/�L#�� ���h��4�kØ�7���r�fk~Ƞ�E�,��^�}��Q�,[Vա�� A��D�M�!l��WW��J�b���]E���݇Ұ?���ޔe�|��������\e������7� �w�H�آ�J@����'��5�)nk "�D��^�)�|3zOhP��^��	)1���UQJ�4Wv���R�hT��/4\cavRw�f-��."ѰJv삈I5h�υb�c_�җ�����I7�pC�\X0j
\G���?���"]�y�oa~&���H�>��tɥ���fz��}�J���+m�����yo�F�>�g�����:ӭn� .8�n@�ewd0��E&b��9�ew;´�[��
���Pώ�z�-��c�y�v�q|�<,�A��xǄT�SC��W~�p���O�_r@iD_�6Qݻ�s��\u��<R�k�Է'23l�Rg��.zę閯ݟ�C��WJD*�#7e�Z�̂���~��9�x�$���7��<�9�?���T�A�~���wxWi�:q7>]cـb��8~q����X�X���W̭���l�s;��h��y��r*f�|��z����;o�ܰ��sx�)ylԁY"����������$5y5l�I��|�3�)��23Fm	LS��ưL�QZI������_|Af�g�W�+CIU�QXq����vU�S@$~�ӞA&<���T��fM���YwK�Qb�m̱���T�a���*�#�ى��F�I ]�̀  �� @��)1���[�.�c��!��ڊ��kK�aT�`��QEp?H�lJ��j����!�W���if���ϥW����;ߺ?9�/u纽ci�ފU.-/�
+V9\��+V;���'�X՗����o�v�P�oHƀ��싸�}x=n4���x*�4�����}�mu�E�b�*�&/v��@͙�+
Ɇe���Z����g1�E�gXA�F��D�<�'�����u�G}w���)�Y<������t�#���_qQ&�t�b�U���**��J/�~�f��6��D�u�0�L�M�)����n\��N�im��4����U�O��{���(��J��!q|��z�H}.�D�DI�s�o�g���Q��X-id��2�<n�[��/�a�f�XmF�6F���C� ) 0��	k*��}�������e�|.�������͡�OOzʣҿ������Ng�ufa�Ԥ�u�a�_ȼ��p�IG�z^?~�����/�R�PF5>plԑ��Dn��TS���Iċ��Qu�����d�����}#3��p0� ��A����shb�b�1�4�ޱS�!�L�Cǘ�'2X�75�:6un����uT�E��;*�|~�0]}���}�.���X��Υ���i��?-�3#u����q���6N�=c��:˵�.�N����f�Fu��'{�h�ޮ:��D�`��+�v����國sW�<@�8�0b�)`k�M��vp���ͺ@#ܭ`aVW�	���_e���fL�!�s��@o[�_T����iFs��������˳s�t�Ż�Y�^�n���L�qSg&ϙ6*�n��y-���R��0�=��O��C�����Pb��sLc���8�Ք�ԙ�;��6��&��W���y�Z��E�q@����m���F�v���0��i/z����+�t���ID7�>Fk����/f�ѱ��7����Y��q7�9\��E� ��� δ���}���T�$:gG�����A������-}�;�����M3s��޻���eί���/����ԊZ��@�iQ���+����K{�n4.x\`������������4p����:�Ό��.m���ν�U_��A2�Q��	��L�f#�dmH� ����Ju����m.c��8,�kFC]TM߀6b���y��3��D��k^߼��t�_|=�gKY�Ngwcj8��Rf/--Ri��:YR����fSM�S�+=����ځ8��~d�yғ�Tp�M�d`�Ȍ���Ȳ������r�ʪR��$��Ҋ�B 	#$�	!�1k;lf�D���3቙��n�{"�1�&�=xŋڣ��2b�X�&�RH�U�de���߹����n��r�L$���Ro��9��?��1�DԲ�1A��zL��Jrw-�asc��T��v4�[et��)1,�D`�+�ޢ�۽`�{��Ŏ�������Wy����L@���F�dI(�tg��}��Q�#����
�ӟ�L{��L��¿�@�8��}���h����/3w�Y;rx�*���E�;��7��Zb�]���s��(5����yc�6!��� ��Vmh���ă�V�B�K o.���}��7v]S�y,iF��3G�$(.��LR��浤DU�`�(E*�6��������w��W���wJ����pkAj\�}���K����LP���-��_ ����	ϡ���ȋI��趕3Yx@pUL�����?�~#��/�R��ؐ��y�5�p#E���g�
0��_G�)���ø"���F�cUdֻ&�u�N��N�2<�Z��؅0������;Pc��i�3qxϮ)[�De�(�D&U��N�k!�q=�0�J��@�
��#��2����[>��:'¦�C�?��V �r��ӧ���O�f�`�Y�\	s\����K��f�5�d�^?�@=HϹ�+��_�^��u�RE��T��4��ȧ�	ӭy�C��km(\
D=��m��@�����,��Ԥ����"� #n?��|�"���"�6�÷��.���3sԢ�N;�jVo��|���frpWm���|�*�}aN�D{K7���+�^��\W�\��j#a�������g��0b66��J��ؾ�D<�P������g��+:��W�͠7���8���ګ#"��$fg���ِ�'�z)B��'í�!�K���L�Ag��@���X�M^I/X��r7RzLO���&� �$@��85�OڲU�jV_���#ǭ:1c�V�z��v��@�2�IA��D��p�C�\�QQ���8J<��_K��:��ꈥ����leD�����d�S��S��B��Q�{��ET/���6�ݻ0-#� ��}bڎ?a����rXS��%o�	��'S(�j��i�c���*:��a�b~��T?ZK��BlvHҤ��qc�C��y\�{�H��s �T���O�6�|<W=��
�ЩY60�sQ��N��k,��(ّ�XE~u�
t�F3�`���X�Y]�^�Ʌ���|gO�-'v"j���:�!��e/pK�u�7K�L��'���UJa'���!ڝ��}�f6��Õ�9;���?��#�:\m>E �6��>J_��+�����J��L�Z3^�/0՟���|//-��x� ��Bja�.�>�l�Y8%��|���eo?�n��%v���5�#z� �Y�I�)
@'P� v#��<Y�|`�����/��{�Tr�
9 U(2�-!0|�Y
���RܗvQU��<P�XC����W֨v�$�^���I{:�r���ZqY1B"Z��>�������_�'q��\�zΐ��@�K���޲\B޻ m��@����]��a�hu欓�;x�����_{o��ɤƦ0�[Mc}�,:h5$jM$����������a����К�R	m ���rΫ�._�����z��h��>�e܉�O[��`�j�6o�loy�+�U��>��k3��T�@��Y��rS~r�z+%�2f��e��sA���u��l��7�
����=@����x�8"��:Nc��2/D�����*�ʟ�&F(��,�m�\o�s�O �Nf��Z�bZN�t�dgR�W����A��%��x�(�׏ϸ��`�Y����Oy�=�'Æ7|��1	b�FY�];��J�c�d�S[�f3�n���[��軒Յ.{#�!Gq1�!|���a!?^�"����(�96h<�~	x�3�j5��rA���m�<k5�X�����42����~K�[l߾zn �t��@_c�&�����20{젚��^T��� �0	���SQ	�U=t�✹&@�Ď�^AJ�i]�������~
�N'�\��70�-��kWzX�ۄd`P#�������yp�� RM����T%x���lI�A��B�n������l�[n�:습���v���WZ��l�&vx5���݇��Q�<?��w��Q4�h��9y��=s�{�]��=AF%��ǺQJ��0�[aݶ�6Q��q�ngE�x����W��]q�Kl�maΕ�L� uv[�Z.j>�G��(�P̛����9W�DEo�(F[ ���q�W�e,S�>����6Y�`/�&]7l���p����jt����A��~/ZD�����-��	<|��>�Ĉa�P�E�����}Z���[��'�x���w�զ'7[�r4�6�<l9��WJE� M4���\�0���?�/��V<�sL�gi�Ӧx*�ޜ�?�Mb9 X��d{3"�z��A��Bs{�d�)��v5��i�����J��r����ޯ��/�gs���_�2H��1�p30s��Mo��n����&)�3!^U�DEb"���H/=��5ߕU���1�:����=��/�^�#!�ƒ�-2�Ҟx���GK��r>�8A�*�����Jr����b`� �{
�}���&s<�[�m[w�S=i��������ο��p�J�̇�N���CE.�G�y#���'�7��P1<�/B����s��h��o�ɴ�EYW�zf�(�X ���"������e2es-�]T��̘� `��>��v`���n='���/b��S]R6�����^۽߭�Z�&5�"D闯�&WL�_ᑷ5q�2���^Hܸ���=�y�s7�k�.U�>މ7��jJ$�7�sG~��8�;�{=�����Hw�c*��E]�o�~ǿ�ı�yX2e�����_&I5`������ӵ~ވ�j��J���@9��I��z�i�������$�C1��O�q��j�<W/	�or�7�&��U��B/���@�Y�7h�o��"�� .h�X�_t_������'҂�����W�)�iX��\fv�ZSv]�*Q�011�3X��^hԛ��Oe* �YX��ʞ�d��_�
@��4wG1"а�?����������=��Q9Y�U1��I~2�z�Bq-���������/��}8퉙8�ʕ�.��۹k{xo��t��V�~}9��"�<�]�[�=��O~qkg����{ ��{Bxg-t/�d��-N�a�i?a�!Ë�:��j)��_ۻ�s�ħ�/�G?���`T�t���W1^��g染�,λ#zfE��v����E���Q7�'a��}�;��Fy��/8���^��:1��j�
�����[�;�EXj�+���Qs�8��ڄ<���or�I����,pdE.�����Z�IEU������{&�ũ=}�i;}�6{�O���\p���(���u%�ig�o���2�[��" V[��P��s�꓀ƃ��"�i<}ٖa��Un�=��Kaq��f��C�ߨ��B��p����"��9�9�^>�gy��1}���W�U{�$��o vo��QHs�?{?��}nkKX�[1,���6��6��j?��[��~hG�խ�:fI�a�f%��$�eU����W��=ޟ7L�YOZ�\�߰�S��r�=jw�R�k��5�c�up�����;��sv�%[�y/8;L��(&MLe��-���p�J��(2���U\�9��yqT���X/���_��׵�3�F3��},r��V5>BI�F��g
�;/m	��o��R'���6z�H/�K��P ��`��I��W�����"�΢$�LR��jiZ�� '� 5�L���y��߿~������y{Ίf�y�! �i� ���)�Zq�x�f�r�.5Ǉm��1�QHcA��rF2��-�P�IQ��5���S�m�z?Q�����v�i��~��sΌ9�X�[���U�����Y;v4tvi,	�X����٢�������@�"Ǩ1й�ĮS�D�g���^>ۛ^���{q3� z^-N�Q.I�|tm���;���{�aݛ�DG������˟�!xc�f��]	g��� u�R�)SB��n\/�2��Пٖ ƍ�V�{ٕvڶ���ө9J�g#�q�,J��d�5���Z\�K6���AK�?�v���%#�hʸc��R��*Z�}���P���z}�?����そ-�,J��a�}�DԋA�*ۉO�7��7�f�UȎ��r|M��e'�fƾ=ŅU����1g4+��8*n
zv��w��O��^* q��+��7ho����?k]S����(��{5Ű>�;Iҵ�;IR#�;^}��QR��&�$!���VQa~�VL_����[�,��=��>�����֌I�[��"�N��ju�QNia!l�]���������_��r�Z���.ُt0��r�=��T<]!��NfolO$~�{����b'�J��|������|��B\U�J$C9f��sv`5��Rn�"�S���}<�P�,+��Pa��E����K_����}���A��V䊼�<g\��.W�T_4��,j�{�N.WV*ZI�>
|�a�f�5���>A")r�(ɍ�L�GD��z8��TT�����&�K��J���I4(�����s?r��ү� Ҫ���)t�k���A��aR]�y?Ӫ�����X���i�gp��⮏؇>�ak��Z�bڦ�7�UW���\p�5[��)�5�>�w�D�a�����U��8�Y1LE��4�+�%G +�b�_2y��{Y��QT}�W/����@�pjo���!����ჶ0Oٓ�0qjv����z��l��C��o^I �e�n��D��$�E}��d���s���< �L��b�J�_��m����< �"� P ��r����W���=�^ �$D� ��|~��⺤?����??r�@�������ƈ���8s�~ ��e�+�\� K}�Ky����RO �ܟc g�!<�M�~��D���򒍣����D���&lQ�09U�Ns��	\/Z̪5IY�mZ����=}��0U*fn<ƭ�s�Ԧ�S3n�8R���o� �MP�N��J(]%j��	N8)����pd]O��"�V%d/�	KnT��0�8e���l� Z�<���x�x p#*�B�#�|)}�>H�H�I�3�Q(Iw�1 �<����v�B�bY� �!���$} �'�61�C�u�^K� �~��u���.5цqEu�(Ւ6C�K^���o�̓��92'8_9 ������w�7%�`���"�2/�@"���k"��]f��}+�������L0�h#��h#���+���6����?ǒ��{r,� �	k�{2wi3k��Tƞ́$2 k�q�����_�r{
������w|j4~����uJ��a�F7ϰ�5լ�ZxtSd��j��kA
	��MQ�#KE���'�c"��j�y5�E����E~���}}���>� �+U$�}�+l���)V��><#ի��t��X�u;��p,;==K�3Q�<I�(&��_n�^zi��|k��`�3AI/�����n׿�;"xS��s�+��"r=>�`�Dz@��E/z�IA�J�mǎ�0��m��CN�(�M�O����7��3�ѵ~*˥��W��O�FLyOx=����|_�qC�TE@/�CWCE���g
�3��c����U�u�ߜ�Q�X�w1��1?�r`�q?�x����[����7P����CF=y+(_,m%/�R�z��P�[ 5�q]@S��5�Us���b� �!�2����e�P��,�	��)R�E����l�36���X�h"�&lێ-��+/����\km�=�0��Jo̕��3	��gI��T�����͑�����G�#�LT���K6=*� }�I{���:TL��Vj3~�G��E��讽N�RIڝ�M���'����n��^xQ �kbZ80�k�d�<&���&zB�DDB&c��B�g�g#�������}Q�p�7F �a ��\�EḰ�� <Q��^����D%�Ī��Q%��������3����
���Im��~�?���N�YXԅ�[�i�86J�Q<�$=x��]!�S�aj&�=�L���	�c�Ј�,0/��V��H t�|f����8�9(�8�y�F�25�#��1��X��E*#�a��\-t����VF/Iq�Q���y�C<�r�;�t��}���Q��aé�r���2��܉#�%aOڵ];�����F��/��Z���0��Mx�V�Z�6=#�2�[����I��V�4&��+^�
���ۣ�8�ӗ���1/0e��z��C������|��:,���4���x���Y�<�����v��),a��M�,�Ns�n>�l^t��t��ag:�W�
΀�!�p`�Ʌ�]���j�}�����ʎ��"c����Q��w�i?��?o�''+��u��H�-��h�����ݴ�w�<,���/>m�f��E�jŹ�>�F=p�)���֫5�u�^U�d4!5h����NznΨ�5�����,nE���s�3��� ̢�w�ׇ"�|q&޸��<wDI�f��X�,�é>`�����.d^�^|Fg�x����u��F_�I��SqJ�bh �J��A�h?��E����0�6m� �\�)��?sԵٙ �NV���F�c�[&�3�Zu"H*iۦj����M+U��Z��e`�ݾ;$�P�UkC���������+_���9�o|�#C���I�>��&ȳG�T��넥�{�,��!�0�G ��Z)�px�k�	��(6��M�͛���l�� ؝��yf���	�>ɧ�I�?X{:���.�"���R u�kq>0"����ܱv1_tO�$��7t9G�Өpן��sׄ���l��M��Hy�p�q�y�r"�[=��N��0#����H-�QRzMMl�V�<�Oj�0���a@�O�(�PŰk��7@���b��es�).�k�P9��ec���9ǵ8���5�
��\����yϢ��zp���,\��p�p�������%��}�o='����0�5N~��S�	j4�1Z7m���
���4�ԷT����߶˞s��>繡�%�Q�+�$�����_�U�!�C����s�p�s��%%�o��Jq<c+@FR�馛�3a��5�^�%FI�<�c޾�/������/�g(}�����%��������&���9�X�ͯ?d���ý^�`Lnu��G�k��6.�,nC��{<�������|�#��?��?�7����Ap�StA�`�]����:e��_~�����oٿ��_�߷r���|4ט(���4L� @�B,�|�m�5�G��a<�4P7�:r	[�3�rh�J��\@J�x� ��yϕ�����g�J���E`�$��F��@��a� �Ap�0��o�}��ĸs���}U�$�F	�̱0J 8�7��b��pq\��dh�I�+ΐ�2��8�L*>֟�����$L"�N�n�#�Gn�F����������{���j�˿��&'�m���"��������$�Vyn��u��W��mx����'���}�8Tm�b�Ĥ��c�d^������u��'H�K�bs��{����VXop�k�����Q��������"b�1�i�2�h��XJ�"]��3vFO��f��Q���ɋ�C�̄G��7��w<����"��t�ϖ��M�y�t���#v�'ﵟ|�+���P9n*����fä�M�Vޏ뽎S�n-4�>7,���=�z�azY��E ^Kf8ԟ$�le�l�SD<t��@%zz�"�1�Ƙ,��A�����\��z衞�!b��ay!��l	�7��g�T 9��& * G���Gnm*���K��fA������c��J�����s���稛�Ƶ��n+z�;ٸ;ڱO}�s�������4+'�Y���l�1�5b����?��`l��/��^��WG	��t�a�P�s�=��s57 l �b~@|���֐rxh��yހ�7�7U��P����a�	H�ؑy2LT'�.�{�!��3���#��YF&;��/t�I̎�N�D�a` �{����4zd:����_��x.��E��̊�;>�x�ĂQ(v�DÞzr�]tɥF��VNx2���Rf�[f�r��񐨥�#ø�a���)�P�/��$2�3�@~���R�9 ��� Wɜ�h"j	���3��׼xj�h5�2h�!	�4�>_5s�{���7�q�=��I�r���K�"-|��w|���*�#��!{�|���q��~��:>P�$�>E2�J�)1?6����$fJK����
���u�)�I�կ��??/�O�������8Ό��-�_lzR�ȷXz[ ��Fg�f���o0~y5�X�3|V�E�2w��
a�k�	'�r�M��	�X�t+t�"�GG�k�B)�(�Cް^'H(����u������-�qD8�l�z
0���s�uH���=�)����6�NY)�����n{.:7�T��V�\�ʢ��tn.�D=��* ����`H��wYS;�G��-F���������~�^�Q�;�"�2X�T= �`?�R%� MZ�s�������@T�u����	�5�l�"����B  u��@�W��j-x ѫ���ŤDޯU�О��5�s뙣0��N��ȅ0|[� �i&�����OX'��|c. ��L[XC�6y��ܐ��m���*�:yI<I�P�T$�1��JqTr��v#y��j����ل����J���	C�i���k��хl��YR��N�T4��Kc�2h�J8!������G���:�� j�c��B k�ypF�R+�F��sv؏���p�r����=�U�������D7j{1�b�������yė@g�ܚ���3+�L�mY)yN��?f��kMî9N
�������N�F�v�bëE`�����^y�=���F�4;|�`�/��.���S���0��,��#�/���XI8Tc�(�$oFa��d�+[æ�C}�6�  ��IDAT�{�jS�����ݼ_N8 �8t9���[e�G2����h�XVj-h݂�ᢆn��[o��	_��1�NZ�F,�.�M�Atmj�do����=n�+_p�M̴�Qϸ�Nhnti�p�#R��'��9*m�E�ٝ%���!�sJ�@U . �$V���=j\�3��Î�z����\�z�0�|Q
7�0����n�C"��+i�!\J�����_�cs�;v��^h_r�=��&gg�n"��U��\�U?��i���} �ԋ0(��N~�#�$8�G��! �^]���$n��:FҔ�^��Ͷ·N��ˣ%�m�5�Һ��G�����@ ��7s����� P@����G��N�k�1�<<)=4�HK��\���E�{l.j��]��l�.6�#v����n��a�L����yu��&�KDU�5�"?Y�ּ�B",˫d��s5 ���Z�"�֥���~����b؞
��u�Q��b��:ܵ%|�����a=LN����a������mێ�;�[ϳ�~�` ް��Sf�w�.y��֩�\�ۆХÄ��o��0���>�v�0e��B>�M82�z�(5�����z�a����n�[.-.�xB��&β�A]�:#�_�ThpQ����������K��p��{�[�b����i��{���g��6�t;�|?���|�R;�[��������a��)|��N�D��FgI#l�$@+���Pz?/�+��(�k\��B���*ǩ��Ѩ�4��1~W���{H��c~��+w��p���@�dڴ90@Uk.�b����}���Y����?�J�6���ێ�B��wZRg���|��	k��s< X��{���{��8E4�ە@@�A.i�� o�	�e��Ƒ��K�Nw��5J�v*=G\i���v��¾3ޥH@Z�pQ��nG�uL�k����aN�~Ǻ�կ~5�������Q�|�3���ǃpֿn����_�;v䐕*d|j9|�m9�:s����Ls�\��H(��,�Ч��n\㢉(5�al���Y>�D���E��ն� <
�W�E�jQ�����b.~�/�� U��%e[�_�|�c������8d��MdJ�b7��j��Tmr*��0g۪��/V�2^r3U�� F\$����ߏyq��-�H�X�!�&x�Q_�ˋiz�K�R22ڥ,o���I��n�V��XQy#�h"��:�E����x7o$�3.':ݢ1�Dˑ�G�O�/L�b���3(ɱ�J}PKc�σ�f�-V�$a"a<(��<��Ӯ�a���9g\BU����ë �,�q��ǥ/�q� %#�Oj����J��aTԉS?�>+1>���j�.v9���j��6�g'�B� NNLe��e�I\A��R5��n�gm����|�N�~��̐U�eR^bY�BI�a���d��F+\�X����C���M .�_p��3C�Ǎ���KF���q������{��R��5�Nڕ�#�����p�sϏb�	�%=O��_��1*@C9\��A�NGu�)K��irD̡�G�Agg$���g�:I���V^?]�K�-P�_��j�H�X��Z����J �ސF���ؤ�ܘ�Ae�řӉj�h��o~�+��-�������)�J�s�Ji�Jf�x����(z���&�Fcr`���F e�%Ҙ����T��~������%i7�7�W��>�ASSS�Q#X�w±pɄ����������~�5a�̎���XT��{W@��9C� �|0Hђ��y��-�(�BZ�M<n<55w"�.����H�� ��=ј�n��%�����̎�O1���:��D�d�#a@��1�	���5n+<��ﾻ��ɷ�{pm�����p�u�f�b��J9��ɔ�����M��C�	�K��W�f%��C"���;��+TG��{*r�Ec�8�wW�T[ƵkԹ�8�����h�x=A�_"�&��e��d�sRH�KO�6��8�G�ݳ1�?W+p��#>}�v�/��?�Z�;�
��l�MK���=�	n��{���Ђ?��?s�p�hH�G�-; �8��+�/8�ڒ�?
��:St�sA"������6���^�F�N��ֆ�$�s��2cO�����^���Fu�SO����>���a���� H �`��JN�Ί~"<��?��?�����ꝏ[�|#dD<�8!];&�ڊUx5�r+�؇��]ĕ� �͘O�r-���������~4�C1N~`t���a���n�=[���V �e�6{�Ͻ�~��o��Z �:�Y�&�a}&��%������E����N�5��;�w3�E-b XA�ɢF�@����%&��j'�va��سgO�d�/� |P�����R���3DFGp��Db�i��^-�	�I�XF��$��:���c�Չ^M7���h,�T�'�T�$r�:y�]��^٬C���[b;%NhW�@��A�c٦&7��][�J;2�ɠ�8�<� .��Vb��aI)��6h�����T�42@m۾c��s޶�VH_9���w����o�s�6Mo�)/QS�N�*62N˾��pq� . ���uWK�T�J�$��WG��^�
��ʵ�����w��3�( ��b�b�Pn�bދ��r"�25��dL�sքƱ���_���z��#Gˀ�FB����B
��X�6�T.��蠀����t�ܓ�Jގ�T��+]��q醉�==k؁��ؾ�����fw���љЯ���m�����a�V�Ֆ���O��A�σ��4�ymCkY�q�&����ڷ��d`��
�q]S�sj����/ ��>S� ��T�p�bʊ�%U�����6@ޣ�p/WO��&Q ��6�?���PR�3,�'V	K����Vo.D�����"G���N�)3(
�``v+v!�F�w�*�Ă��ك���׼�78��2@�Oj�z>�ם��Ժ�m�|�}꣟��O�#?x�����ض�;�`i���M�;��,����l���$��X�� �Z���\îҲ�����7��v�������v���ע��4�b�����Ի�*��u�]9R���J��J����� ļ�������B�;`^!��Yد����Ғ �@�)2��-���H�tsp��P\�"�a��v���9%�� H^9�F��
�O�B ���Q^ �{����6��'�x��򃟴׽�v��=-�GIE8�wx���E� ޠ���D�i*�&ʹ���0>��O��s69qF��b�2x��,�� �:�0惫�//@���4�0�!�D;>�I*	�����&�
?1�ΐ�׆��5�R).��h<�Ԋ�^�8.��U;�>3�Ocu �Vɪ���3�C���2(��b�xQl+����������@. UjA�, JVI��g�*z@���R���V���{roVl�����ٌ	���;Q��A���r���ј��Z��o��������c�nٹ�LS�=�q��R|��ԕ+�{H�VjD�2�B��T`�7��W^	~$|.j>s=��Sp�H��ʹ�
�����.��}n�4��>.u@�\NN,�̦�x��b'f���є�V:9�= [t�@� aY�"qB�t\�xK�C�1��AɿP)� �W�|�'�*�z���|Ĭ6�Yi؅�m;N�l�S��ޯ���)��ōN;����ڠ]DE\cYǋM@2 �T%��-v����_�o�*�^�lW��B��^�1[=&/̏-���*F�J���>�X�J �+^�n�a�|ДWcB*X!X�}r��֞NZ�4�#r�t�U�([ϐ7�@�H�G�x7�������XY6�ex|>
��j������O4��w��t������ُ��z��2ʦ���9�T�F�{��h�c��Sk�:t�<�6��r�>����҉k��X*}^4Lx������#�8����+�Sc���}���?�$-?��w\π?6sIMJE꟭o��->E���[|��L_�NJsHY�._��V{�<�k�0��}r%1!�̫V����*�ʡ 	Q^GR���)l]��x`Z��گs��y�c��� ���o���ਕ���ݑ��LD״ޜL��R�+��杘6�&�<��Q�����1�L ��>�s��Џ�;>Y�`�Rߓ���G9����,��8�-�[@��V� ��xw�!4�p�/;a�N���[�KΰK/=�&�Kv���3S5�cXr߻�%����DrX��F�o-7I��W@L�ߚl���&���姩��r��Z#_j��=�H|���r q���ʷ[�ڐ6I?*䟵 �K>Z��_R�(O�����;��RV�%SH�.}cqS���}qU��6IH̊6X�]I�z>>$]�D�/%5��R����7�{����͛lbj2���\w����
{������3b�#\:kթ�����w�����*Z�&T����
q?��m_iE�C�'�(MWǍ�>�����/山��a	b��<�����	9�m��l��Y|�v��������9�7��2CC�'�.�W[.YV[��J��>���X���.U����xx�b��B�X!��6Gq�R'	�]+$T\�mD ��8�︎rp=y���(N�K;j���|�ө��F_�Sz?-lq��bf.�y�bD�U�C��,����$�{��Ӹ*����K�.���a��E��j�/4cy���b��n�풋ϳ�]fss-k�� Y�H���kw���h�h�9��43��+!yRx�P��J��an�9�F��	�;&{�Cn�}����K����&�v2-�QC�������M��i�Z���>:g[gϲ��<1��sP�#N�W� �}�-V��L�,�Sq�J$.S��D@ ��X�ճD��-p����%���(#վw�����H�Tj3��i��y�R�S-7�kN���j���ࢴ8���(Jn}�(4����^��D�}���o�z�r���m0^#�Z�**È��#���FO�jeҞ�7g_{��<�0�l��B7[703��1��Z����3�Tb<����o��Wh� �dFp�˹�l[?�[A��Q;��Z���RWxqP �wT$5�|�.ngs'�W��v�:h� Tu���g�D�F�'7e�"ba�NLa�Df8/���*	)����������1Y<�Q
Pe'�q��	I|g!(���ŕK� (��W�G "}1�䪦"qO�*ݭ6��A{U ק����p=�)�c�VMqഏkpm~�]��~�-\[ܳ'�M`��Xc+���zR�����1��6L���b(�����p�R6�N��@Kܼ�U̢�^�g�ev�;z���߹�����4�Sj�I;|���}���u7��]gY�4��b<Ƣ�/�8�� ��y߼$뙸�H:����\n�9�xUߊ��'��������M���vs�Њ"?f����>wb��'�:Ĩ01�h���	 ^�n���s������	[?��~� 	���cq�X &�^��^�X�8� *�-w 
�)~�J~����$�^zit�Q�@��K!^/������x~���8�w��{"�����M���{|�rJ۩���'ek�$��]ʅ�爣�t�RPEW�� �#��O��v��2(������n�#��$ƕ��MQ�p1�2���H��u�;!���>JGK�i�*�r�+��N�6	t"��"�h3�*T�gGpנ���2^�햔óճ���I�6�FN��X��^I�U��'m ���{yھ��w�G�.xS�Y�ͨ#�:�#q�^�(R�.?�8�w�%^�9�	\�{�����5��sZn��%�T������u\6�S�5�-kwI��-��0��NసVu*��rFT�]�I�"���ʑJ%j���ű�	�Q��N
P�  ����>�� G\v�����ߜOi�����+��"�/`��v���  ~�>�`�� m!3ɺ �.� Ĺ��`M`��T��K{9�� � �r_Tuc�����f��崝1�ܛό# ��*}.?S� ���r-��f��f$� �6����@9�񑏻���w υsy�<��&b�1�;�:���z�$��� @�b�3�����G����9�TX.%�N��2F-�AR�&Y��tлD�J�3ʯz��焇q�ˡnw��	Ot:�ҞRO��*�x�b����E�U{u�#Y�ДA�u�]�n#N���;t`�@����dح��a�΍p�ˢ�?�<�_�D���Ćdܒ�	�L�Z�3�� �D�X�$,\@���x�c��NΉ�R% . ��� h�� `D;��-�K,.�������m��s.`�m�x��q-H�5zv�E�JWʸ�+���u�I;��6p]ڦ�d�4 j���6 `l!�9%cýd�U\3@�̹\������fD{�� ��OWc���<S�XQ(�TO�������`֓�;b�S5k�p�u�<S��;�0*ktӆ�_��g�c�\}����9���uV�R��D_;�	R�TORE%�Ai��ԁ^R�h�@��ƌ�n�B�wB�b*���muc"5���kAIg'qKzE�(�1�<�(~ �u�� H`��`��y\������9'��J%�햛�cS��z��&j%k5J��ɖ���;��G�Y+��="�Mn���W@�� ��{,�0u�҆�Dn?�;:�K�'�����쾺3�	��BC!�ø3�(s@���9�c/�<+�hh�D%��$��Y�� ����/s�Ϝ�=�N� J��xp> H[�tʊ����q�@��sƐ�܇y�J�|T2���U���O�c�#��VF;qb|��*1���޵�����C� 6>�'����G�.���).	s�����ǣv���so�I{�-W��dhC�n��R�[lrb�-,�y&���	c���G%F�A�#	W�S����|�Oگ�. �������9j�C",��]�*�{ch�9�n))U˕�g9 �lpR,�t���*E�%݊&��E���a�8Y����t�,UP�N��]�;`{�O�=I���~�v۱}6֜�v�V�۬�[���1��s�>aϏ&�����A��Ȋ�o�	q�qg�XIO�o�	 �ɨx{�ѽ!D28�y ��3D)U�P2����K[�r�&��ui��^����W�'O�B�űÙ�8SUX��T9^_�O�6-T&������㽌\���r	 �pќ#��r�p>=���4��kr,��o~����I{�'����b#�06����H9O�gq�P!�v]�)��UJ�5�l��	��bpu�[8f�v��O�N�ԯ�����a���\���V�6D��v�|e���@ء�^̋���xx?t�����P�Yv	��}�Oi�������N�'��.��J��KY�Z�U�?��N��w�]�	�B�=��.���jb�kP09`Y�e ����鑊�vSQ����!;��vÍ�И�a�[�Ul~�p���p�eu�'�·*�_�\�
�3�f�͸*��W�B� ~��+_g<�^g��H���4�p,|~c�s�V��3���(��Z�<x�'�����N\���k�����f�zCB\�<+Tq�X��Q &�����9G�>��NT0R�p�Bh[��8��~P�	`�g�ϱ�j,�K����5.�˜��8*�>�y�kȅϯ�����c��-�a�զ�9n�G�m��?f���vɥׄ��u��Zb�z7��"�$ϙ��|7�օ�Ah���}��T\�gc��O�m�k2y6��4/�!K��p%�N�ֺ�r�SI��ݥ��%I2	M��o?=r  �V�5$�*�c�9�ゃ�k����K,�$�L��0&?�0]��2�(Z�����q-���B���"7�o�-a��ڑ�lfS)<�N�QˀXE=#wrP^? �����&���r�J�˱��G8+���� ��=L*��x&;�	�p<�l���\ �de|y��$�ȆH)��\�x�<s 
�gŽ8O�)8y%a�E{T6_ �v�0����617��ע��ƫjJ���C�i�Wp���h<���W�1��1�<��8T�)�8c+uc�x�,�+m�m|��d�L��T%��gB��ӆ!O�u���~��b�l�X�1�O��b�>����w���֨W�~����v��o����R�<���`�~�T@�� ~�y�KV�"���j<4��K��ld|׫M��y��F��#�e�+r��Zµn'�R�s	�!p����v�,����.�k����)�� ��o�ǔ�c�P���cLbb2�$���K�����U��7p����8pЧ?��\^"�(gu�	�,%��v+�;����vϧ?o�yͭ1�O�Ӵ�MC���:�����[��0F,x9������?�X�Ð�X��])�����(%�:��s#LD&(�v ,�ǳи�:
�г���t˼�N�$��㸮T
����C�^q����7��g@�k�l ���o��y1�|/� s��.��`^z��IZ�pO�Oq��2�%�}%Y�_��I��gmb���U�z�}qf��/~�0s�fd/(��u��U�am���S�Q��ԩ/�����=�������T�t+'ӱ��f�oe%�� K�qw�qG�����!)in���{�9I�+{�|đ� o0HA/�S� �1e�W�B���=7I�2@��T�+�%]�*�0���Xc.�i�p�<Q�s��+k\p�E�E���!
�O�!:&�@
7C� 
�]D�4�p��	1F�ǽH�|�7Dq�kHL�V̆��g��'�\�&O- FXDO<f\tVh5�8eN[_�����~�H��s&()��p�^���s�3�OARoh2KO�݅(p�2�
|� 4һ�;���>�d\��(	��) 7��k'5��?�%N^��?�M�`�'����"����K���2
�~�W�\����MB���`L7qc
~Иs��q�0���$$�D!��j=�:O�M�x"�#+��j�yZ�	�0s;AWO4�-# �Fla�y�k_�����7���_��h$��<|$����{���o����iH0���#�y��`n�����ճ�z�W����{G��J���R�8���-���XE�`�����tǄ��Q���&5�V�X<tL�*E�l &�o��oG���^�:���?��k���o�Piw*& )�L��τ�|�.��t�𢳣:��l���"��,�{&9ur��J?��:�/����o4Y']�<Ε�����k  �X%��\�+xC�S�%�{�I4=�-�M%��.�N�~s����w��T	>���@��~kj��W�s}��tw��i�)��kjQ���8E ���&�!�u-�Qu�I94��q�&�st��W�K�K�ubn>����NEIy��;m��h[1x�"�����Q6�'�O�^ �+�XA�"� E��Cf|��К�3���*<�Z�瞽!�k=��Q�^������C�k���@���ђ�p���X�ʅL�ո��K���1=��
~�|�m��tϋ_��o��A;:�����>f��[��.��!#�w+iaxn��p��mb*v����{���Mw�y�i�a�3�r�R��rN*���YC���3����E��G��G�����=�h�c�}"�aM�H=����x�s�
�+�&?�ݑ��Z�i��%�(oȟ�=n�ʵ����@)/���,JUޖ��R�/N,��J�����a�z���^���I�T>�k=�����,X��h�R5��nD�6���U��;��}v�ȂMLZ��C{�S�c�Uצ^���h�;��^��F�����_��CG�J��ɥ�'�B� ���1>��&�ׄ{����o�b����jkN0!�ݩ5vQ�&jUk/�^�'C7s�aW`p����bO��B�iBH��$B�HG�%�R�����ϸ�� ;��� � 2���}�}�*��g`b&kv�ۛ��v�%����1`��Y��8���'^p��][���o�I�*���Ӱ�x�����N�c��ŰW��W��ڤW�J�H,�P`Qz�ܠw��QM��}_�F�߆����v�����1)��u=��k��|��~�-������^m�c��J�i+��9��*���I���DVmrz��Aj��*�5/��~��������q��m�\���P����f>c�Fs`^+i�ThzN��jozӛ"|��}��2.�%T��n$)�5��M	]�ʪ�,TZ��X��<`�6g�Q�̑)�I�_�.jI���S��4b�2A�β#��t
�I<7��g+w��,ƀ1��Yq�pw�}w�0����-G��܀��D�����Rb[wL�� }��۱#�6�y{x0-�7�<��-�Z醋f}*�AkA���5^I�R
LWg��������T'��vع{���?�Ή��'�mj:K�Z)�֤��b�@�D
�6*OT� ����ƜB�yEj�0:+镘6y�h��+�א���_hp�{t|&��C�F6�iH��j/� ��l�F�L�ð�J=Ile�؉����DW��Y�pź�@��)b���$���x8Oj����%DN;6ޡ��쑇�N��Ѱv�Px�m����ID]���Jv��nu܆���~��l�=[��z	�p���ѣ���=�����*�n��F:�险 IS����K���"y�H�º7b=���+jL_�G��C�k�pˀ/x!5��aĠ'�D��M�eWP�*�,��̛&�%�n
Lv�P���N��ɸ��������4K3X�(S��qH�|Fe��d�fgH�++�z�w��Q1���g�$B`��J���Ur<�B����lM�7�}��k�a�MTÎ����I3�N���eJ�c��X�z�σlэN�A�l�L�6�@{z��������]�G�o��]`�]���%_>���zLeI>a��T#RN�fP
(Y|/?ie��3�AZ��Y��>��0�'=��G��s��K������S�k��hRD�7���+� ��EQ;R_x_\����^~� ��IB�) �?��?���>�яFu�9�3p�8��.���Mo��`f�q��ܿhS;-��lf�|�zb�3a� �M��i+(m4H=\<�67h����nVA���ٰ~�n��Ԍu��ӭL�x��>N��f��J����XC�h���Ry����3:]�{Yìk�<X>��OE��t�rS�a�����e8�1+H���}B~�5ہq��ڃp��q��[7�F1B�R|\6����Y\ ���y�\A��c{�SH�p+y����z�1�@[ ��N+� {p�|��d �f �2b�Bh�p�.�ռ�\��a�;bm�����\?���ؠg7��\�
k(H�ݬ���d��S���歜�����vn�f�o�7��pl�q��rC������;�c��^��UKF}T������䋷A�;�D�3�	�꣇-�R)|^���J�Y���_�L��Q;Yp��w'����+������z�������=��w�;�K_�R{���B�ey�h��So�;�D���$:jIe��{�b,@��'73��#ùS6�诺�q��қ�Rܰo����mг��:���4�`Ǐ��v�F-s��t�T �ik^�%7<�v��8�i���j�u�}�=k��W��r;`��B
�Cc>^Q>�V���E�D�*I[�
k�y���}��T�]-W�n�j����	�y]�#��V;A�6�w��."���h�"����9�o�v-�E���+�J~����?��N��R�U��ꂼ�dR
��> ��ІFhx��l�&'6�wz����-;xpq]�����'��z�S�ݍz� ���Ӧ�mo{���c���I���Z,��l�lz�Lkf�Ըa%�'��T�eyT�
C�o�u"����3�>�$jSHҲ�	�A���w�ԧ�QT:S��@���D�:I��D�Aة#�IT��J�ȳ�y6�GwIE�� �+6���?�{|������y���}�I��
����$����f�mE�h�j2�w6�9۶���0/)����I�C��½&��J2��RF9=<��
1��J�$�J��g�����S�7�'6h�i��N�Bnz�@$��V'���k���g��/<C�1ĵZU{|�U&f������z�b�F�T�6vDӱ���Cs ����f����������/^c�S�#q��-˭<#8߫E�6�^ .�֟v�̱.qW��y���'�H�Ġ��^�je��8"Kv�
�KΉ:٣O�%��Q����X}�+���s W>+K�t5R���!:#`�w��X��F/��"��8�Z�G�_.��L��#����]x��v�M/�͛C��cG�
�KF�0q�R�3�� ��<n��9o��mp�]��'.bra&�c�R�@6 x��i*��;�T�3�1�J˶l��c'��?�����+��Ѷ���`��-�N[y*����n�lO;mG\D�¬��y���ڽ���ɵM���`��d�)Xs>�]�
��L*<���'�e��e0�Y�$O�ߍZ�Ռ�xN�UNcxa�"�~��N�Z�}AVS��а'�Tt�D����1��j�XDՀ:]��#�b�0a������薆h0)q����.�Ї>sI�d<\��[����8�سx\7|�e�t��G?�����7����s�ґX#�رV>Lr�
��˃����76�c�q`d�/�`�qL �q$��mг�2Õſjd��������~�ؓ���W�������R
@�Uo��a�#7�l��������7�9d�(�>p_#�Ǒ���D�:�%%Q���8c�8�R�zݰ�Q�(>�s� �rM/�gx��:�j�Z�]�3@(ƥ� 湏�m^|Af ܇���H���dm��ݞ�:;~~������H�z��*�΀������_�r�.�|�!���@Qe^��-ڎ��؁}���){�˯��\zA��ь��F�����
g���p�
���:�Z�X*�����J��#@�C�E�|�7h�~���`�K�G��0�N��'���}�{�lv���P<���Z��zc>O�s6x��|H��k��62kw����R�]|�����-�t 1O1�Д'VH�7�+Me1�;8'M� ^Z*i�h���#hI�tC���F�ވ�����Ύ�,��*�*��C���w ��?��_(���J� �<j���/�F9v>���^�̫2�y�4�_��6w��Ϻ:؈���'��l��4��G�%y}�n:�М�!���f�9}�}�} 6}#��6�ڠg%�[J�i��k������m��>�P�yr&`C3p���pV)i���a}0�J��}��G׶V+� w�_%��^SPG���I�4��aV�I��UN���7��0�!�s���+>�Ւ����r�i��t�h-�U+U�(n��&{�UW�J��2���]�݄���p���۫���>��A ��j�](�������$�����I��]aמ��tI)j�;�o�2l�ਢ�s���K=1���sx.��=+�u���Xk.�/ʕĦ��A�<߾�бhWR� �S!X'F�Yw�+�ֲ�Z��r1�E�)g�`>�L�I0j��)Ҁ:�"��{P���8��a�9B��lujvr
�%9a.i�N��I;>�E�5��c��j����HUdP�T7L��n�q
C���|�)= �M���n�\Vy�RL�A�Ӌ����z��J���ѧ�~��]�v�o�˟^l��#sV%�`���k<&��{��MP1�|�
��J��A�l$8�t��r5����t�xo��F{��O��G��l���c�@��ԗi2���jL��QM���y�Y+W]uU/�?��)��d��mF�W1�
�� X�u�W��b`� b�}�.��Ҫ�Q�t���Z�10�1@|���X���5���)��p� 0�p��Q���������NBf�.��}�ԓRT��D�Und��>9U������9gO�UW�g'�"�[�N�����@�j���?ʋ�9~���S2δ_~����.j�LS&�����Z���m�4k�]w�]�ޫ���+��18��LF>}��k\0 
SsG�%�W�<��4�~R���p��L��t��ž��RQp-�
�J	g���>�ǹ���#��+������f1���Pi,�b���Wg ~���j��-�������㚨-H�9SUd՗�o�_��/��m"�`A����j׽�;����N�s'�����7�3 p��FE�� �H�{"��HH.6���£���T+�x��a�7虢��f��5���Vg�R�f��b���>g�ݶy�:Lj�,9)Jq�v"x+D�x}H���d� ���+12
ʐ���WN5��H��6����\e�P����7����S=MW����c�[�� (�c���L��>��z�Ii�=��tU�ŗR	3ދ��<���&�7�#�Xd7Mc1�>�&�K�i�Ҥݲ��ħ��� *��ih��{U�b�!|�ѡo�=[)�}�lwb�j@\��}��
�;1����f��)]�l�rukTE���h̋�[�ը>T)4�-~A�]T�Hă.��u,�[��:xCls�F��0;0���	�� �F�p>�y��=�*m�g�(S�F�(�OI}xG�r2����a�ޱ���y�,�U�6՘=���h�����vp�!�P�
�]�|ʞz�m���I�:c�&
�JqStPlT>e�j�A<x�	�VLH�td�6�YEi)���*�Arl��C���|���g��VZ���g�i�]w��>�b���	�\�ienm�{婴n�qz��Tд�-�I�trV��NO� f�X�A��?����TWk�[Z'��Ϝ��I��48P}�-6\��AyAh�9:��~�Q{�����.�����'�SOcF�Vc1�HFϵu�i�,%�zE={nj�Oe	��>���#�A��*����X,!�A�l���mƥ�5��۠�C�
�����}�o��O��B��n+��ö{����Q�s��:�vO.J��@q��cJR���{H���[#�9�^'�(��D�LAn�(���@�Z��G�)��8`�
����O8���1	��� mҶ�R��� ��N\��.�#���&��q"�X@[U2'>�
ߠz6SVA���$-���CZX���� [f*<�p,?\Ӓdb �Đu:�k[�ֽ�0je^�w^Z�I-*�$���b=�y�X��U��tu��OY'�5��)�2Р����uvyNЋ��|uoo������rG��V_<'����hյZ�w��B�~�Ⱦp,���#Mb�����$��?�+©�'j�zUF��;@z�6�YI��j\X�额q�Vۺ�b��ޚ�s��]v�U����p�R?�"	��Մ������5���$�� AN1j��O���H6]���Tii?a�DH��Zn~ ����V�(h�!XMt��z��v�^�<���޳c6�W_n��-�Ś�j���?|������ر� {)��HO���"�̠rV�5� ڢ����}�7h���T�%��`�mˌ����[n}~`[�a=um��67_�a�Ie&�#N��)=%�����n7�}J\�d�Mѷ����ٽ*B@*ψ�qN *�Yb�|�Ȩ5_���	���#E��:?D�{Pw��� �kt�?z ����s��f�!�e�v������	�N,�Ƈ&M���U��N�/<��\$�`%����ʡ�ngbX���Ǫ�N����x��2ܩ���U�^?��\��jh9��Y��^�u�l�F&�X�`��;��3�w�Xu#m����v�pÚ��=�$>�oV_��,P�aD�K�A��t˒֚����^Y�y5�O
�ϕ﫶g���ѫcAx���C��s�A�+���*�E]Bw�XuZ�Zu�lG9B�+� ����3�]&�U��a�p�jK�d�)�C���m�����+���w�����|�}�O�(�@���rf�����%t2B��B�op�0¦^-�:��I��l�\��˗_�o�*��Q��4��R��R�Y)h��~Jr%��,�۵!�o]�x�R�O${MT�q �g�}N����=ީ�NY���$���nB3˨ۺa�����R;���?����z�.��j۱����5�;rׯ�t��Y�~>a��A�+I���F�x_d����g�<�mO�XOb*{�D��I��ז���XPH�ة~��Y�/�?9xP�}U��X03�Ȫ�N�����rq���\�R7x_[��	臹wr��}�l�鿱���y���+���6=���漕p*��=�W)�}�y%( "@ݿݍ.p��K(�fc��}�y��(�m�O�4�7��Jm��/��;�����c~���,^��k�_c�-�1Cޤ�ڻ�~�ܯ˓�4�O},~�w�G6������W��N�ju"���G��fX�����o���g�]��b;��K��8����X��{���4�Q{b��=0|<��yU�O/�lW�>@��N�my#�h6�F��=7�XHe��j����@����6-�Vd�S�s�
x�,H���ي�-�O�V��(��|�-Λ�����|�^�����ZDZ-�]^��r5F�� ����Z������-�]�{F�|𵨓��pN��o)�Q *p%�����n���9C�4NF'��QB� ��Ԭ��KI|��+�&Jm�s��j�� ���u�sk��F�@x-�%L1=��LZ��i����'?g�~h���E��isI#\)e�M�D������ƶ��n�����o._�] -����yK6�`+�� ܩ�}l,�`)�����ʸP*���`�����a�^Oʥ��2p)�Z��T�c��I��`��*�D-�5�f��܍��\Wk-8�n���y{��OU�uߗ�|Ggx�2��D%0\ts��ߋ�e����w��'����ˌ��7�4�t�t����`��`F����n������Y#%]��t��z� ����D�2y���*�Ν�2����TT$�U+i]��˕ؿ$5K�6Ab�̅/�%����e17Mx���>�J;f���K�r�C�j�+&	ދ���jSM��_���H ��D���-u�z(��6��v��/�ZKlb�j;��bg��۪�vb�8��.8i�9cX�DuD7^�T=JK`��h�\o�r~��p%�㊟ך�{ݜcNY����a�e�Q�l��C��1�x�t	�xO7<��a :f܊�LO��rX#1�	�-*U"`x#w�_�gG���{��X�e�ڭ�u�i���b�F�Ϭ&Ղ|��LNs��KI#�r� g`!�TCT��ҝ���V���?ߊxLǈ������^W\qE�
#O��z�.D������ܞt�Өݍ�a�������'�r{r-�Y����2����Qi��C{������7��]x���X��C��7��K���:Ҥ�c&ʎ��wm� O�!��:��2����NR���.�kb�������� 5I����r��uXZ�b��ü$L�C�_��?�jfړ�FQ��=���_m��/9��^�Z�
�Нw�Ҿ��'챽Ǭޘ�fk޺j����Qc��h��<�Iֶa�z�O0XA`��H��0��
�k�'���A����7]�.�0Z���Du��k�F�J�lg�}v ��ǜ��*�' F%J��).�)L�)�C��Т�1��n��6�����x�w��gϞ���/y�/G�6�j�	��㜤� )Oe�~�m���.;�^��Kl��h�Fh��l��1=/a�|cґ�G����M���G�~Q�Nu��2����+����'+�(/n��A*3$�z�68鰓X���9ߓAx3Nt�3���#(�,
mPK,�6����a�fw����Z��d��"�i�����(id�ն=�ϱ_������7	��lۼ�fǏ�#��k+V�Xb�����P$�*�DMb��.�,F�RH��ɚ+}�c�@���7p
�����$ot��"���0�SS�5VGt:\� ��v�M7�ƞ�Gkr"(!��o*�;�������P5��ߒ�g��뮻b"旼�%��W�"ޗ�R�q��b��~�R��,�O����-��^�[��T���F�h|}9\r���,�c)Z���~�䋤c�b�l���A�������-����v*���>��������Wx]�w���뢟n�����̆y��,� i��(z_�( 0^bj�wۻ�h�O�$'��1�O�Լ��� 9���P¨T�F�w��ٳ9zE|��='���/'�ru��@Y	x�/8B�0$v��/}�KG��e[�� ����_p˔bS Z�ت��涬`��q�0����m�{�����}�=��S���J�̐��ΰ�$աc�(�Q?N:��P���J"�s�=�^���/�rs��2���>�у<!�d{����)�ͻ�~9�V��f�R�ӴV˔�?|�)+_W��Zf��"~�x<0D���6�1/E7mǪ%���K�r_�Iu~�si�K���dƻ~�`�+�8�����t`��~��n��Г$���uJ��-ñ<��#�L���g�G�17�s�OJH����~T�W9��4b��Rq�T׷�h��G��"}2��)�I�[���Cf׬�J�����w�"�|�gon$݁y���3,1l?��'��R`&Y&#��V'�jWVs���;��*a,��G����0�m'����l�D˶��;������<RD+���^�M��z�z�9\)�õ�R79��L���J]�q�6)@ə��ԗ#:�{�qn��U�P�8f՞��X�����ʓW���fl���:��`ɔ[���a{�5W�A ��x��hx��I@'}.`�\��܋_��8����IKW��?�S?��cء0 ���cy0��a�<��|�3C�/�wa�,����w�=����c&����2���aB#� ���{�>a����G~z|�R���Y��1��8�(P��n4��� �Q�
��`���{@8U��r�23���/��[� u��Ja2�ݜ�qaR3�}�n��e�}!��ϯ:�=h�ő�d����'$��t�'���Y�U	�>�po��N}���ə��ONTs	�q�����Tع$*�$jb���[:�|�[��{�id��)�r��$΅X��m}?��	�pȾ���>���h8����;ڶ�:�\{�tû/)=+ 2�06���	�.��(�mw�����k��Q5F�+��2�� 0�l���1Q���Nػ�o���3��y�e[o�˽��^���[qΈ����ΞC�Mn��WLȭ����~$}�~�;*�����q�u���9�~~:�Evm�nZ���ޭ��׉zǩ��x�7�Y��?�A/���׽n�v�����K�
?�^�8�Z`ﭷ�:탹9o`��cp>�{ؐ���
7�|s��*8�O,{�XjG���� ��r3Pzn�|�}~CJ����w\|�nL,�������7�G�%��q�q���"`�2ep���g�Y3��!�9��J��o���1	=����~f��M2WT���J��q6<p�C鯾�t���:�6v�����P��l.�n�A7�[k)[�[7QF���8�=]�p����h����r��zʠUp߭\���y�G��zg��b
S{l:�L��섃�g&���ի��,�O�1}��ۋ�@����u�r��9��m����"5�0;n�`�m��n��c���aTY�)}���D��kw�-����&[l� ����T��׋ 9�4�7��w��&���5��0 �[o��m�\��6�ݥtp�ĵ(ӃS���F7=`����ݕ�3wB���X�N�d�J��Zݏ�M�� 7`����������;�i�F�"�Hl���z9,���T.	��>���旁p �9&����Q�;�nq������4����@t�w��/D�$�(�iYII}f��er^���"]e��`~PU1���y����|B�LRC�h���kl�	'�
d�,�
0�c�-�&���Ғ;HKt����u����v������ݻ���t�=/^9�m�	g�h2]ty�����t�iAZL"o������̛�*W `��g^��l�) w7gyj�/�NR�*�<��@��P��T��!3D~�F�ϚBv`j�޺�1Q1P5P%>�&Xiky��"==VǚŊ�?��פ)2���e.�.=
gBh��X�2UҔkPڽ�NS�?�$?+�^DƵ�z�����u]Ϝ���@|� �VZ��=�I��2�k{i�����d�ʢ��]ߠEX�]#:�׌���*��\r��bV�̒`Ɵ�ɟx9X
����o�?��OA���� ��� 6�͑Z���'hͩ�3�������F{��Z�n+��S�+ƝZ��ˢ1�㼳�q���4D�q���(�VC����x�)�iB�c���(�x�����L�W\�R��ot�,���<Nn�Ml͠����F�&Mz.n��0�|v:�HJ����:�w�r1�k:"D���@7;���C���ܸ����x4q�Y6_g~e�L-:)�a�c�Y��ô�������eS��T�t��j�8�ndǇ��d�� �=��)𬨦P�h�v0��ݛ��o��t���7�������0�qݜ�6\E����X5N����6�������^mV���TL�S�M@�aX�g��J����4��4[+#��Cs)R�eb�k�ήk�B�6�� �:�u���O�{��g�p��X�Re�0F�$��5�\N6kM�r!{ՅM�?���1C�5���x�);��x;e�h�9.���bn�k��֣�!O{2r5~R��f�T�Kf�h놌�C"�����%X�i�$7�$e���&`��,��g0�^{�4u	6~C�����+L�`��` �t��m�:��al��Z�r2��Fo��G�������j5L@�$���ÃE��]�yԱ)p�=��WC�ѝO']Q�0�����`g`�"?`�f�[wh�_۠��R�/��Yh��d7�7��)��� �ڌW�U�&<aM7%(ޘl�&-���U����	�%�w��`Ǌ/f*W�'��@a@�!��+;(�
�^#cR��D`'�\���y��I�Z��ʺI~�2���r!����*���SG�y(_1��?�����o��-�T����y�SGdfХg+r�9('��9󩗳#�	sϵ,-7�l�����^�� �XTה�C��`q� l�L8_C��,�&�ՙe�u%h`e��05��Ɠ\�&����q����&���Ν�Ƭ7�wҀb�_z�F���(�!�Yk���E��/�y ��d:�S��׌�,�M߃�|/U1�ħB��^��ċ�T�Mv1���������X@@��x�K_�{���Nf�	��Wjة{��>jU�~�4 ����f]�E$\�i aDv3d&��sB�$�`�Y1/GuB7���L�z��1-�E6>�'��I��?���/��/�Q�����漊���G���ƄMjV�M��M=F�0v�YXX�L96X���&u�Ė��s�i�S���ߑ	ov�0��]��ls�曞좲�Q��zn�Rf���-:�ڰ�ONIU"���F��0j;��Rׁӯ�0iR�9�7V�:C7�R�Ә�w�^70�pV�{9��N�(;�r��4�����{���^���:�(�iH�s�� U�
�E��`�M� �|Î����V��ͅ�7i"�f4�;�j`�,�,g���,��<S��l[,-�=@��ݘ�h��g7v���|e��'��j��>&����h�NV4�ko��38�βobc.��q���zӨrF\����`ves_u����m�ct��p�MZ�K�A,?E���ϵ%4�����k���{DǍf�F���w���h��3s�����?O�*C�t< �m�N�U}+c1���fl\NS��q�{] \�#��S�z���*[Tl2r���r!Q:�dZPؚ�KD�����U���~�{�s	H��7���Ƙ%86 ���񌎘�9b�p��G;��!���3;�\-��C��iV�`V�=�W�t�y��w�!�`b��k�R���s�Ygo�EY90M�{Ӿ��^�*7�tӷ���t� �y�c.H^t��ڄ����ܕ����w�K�R�������=�
��t�y;�y{v�]����8�ԛB�`�n�)�{�����t`ߡ����vl�k��Ҏ��}�:3��B,AG��rz�����ޞ��=�q��V��9��L�^r���p&�H�)��BsF=���Vc!{�:�9;ܹc)]u�S��h��Y�ày���r����ӏn����ђz��+.K�G��j�QҘ�"�{�k�������<����5��\�']r�cz���MtG�M���O����v�����a����.��ϑ���ݬQT1���V�������}����;۷��'^�ce��j�*�ܾ3�|]�s����[��H�:5D��ID�����[�n�N�',gg�g����{����$&�:�C�ػ19ֳ}�N�\��I���1I���Xh��������+.�Z8#ӧ�a���}z]�|�h~�[�?�=��v�m�m�3vs�� ���MjB���AP�� e��Q^���s�Hm�B�򖷤?��?���w��镯|�w��H͓�Dq��(��у��o���FI��ǋa�J�[����E�xvO3��qV�j�*5�$�9��$�5���`���7�"=�9?al���*ؿ��vdlhh�뎝+&��������?�A��m ��=�)����
�L'��Pڶ��:u�E��qR�x)������ޟ����r�������}B���~K:��mv�5��^�Nfs�%����t�?H��;�o*Lc0�u������ғ�|L�/vlْZ��Y+OVӶ���߹#����?��H�{�X��_v}z�k^h�q6�:���n������O����L+X�k��	�����v�*���t�u'��c�q��*>�_|��?���j ` 5�ϯ�ӿ���O?��K��u _���<��csxם��o���j��v�];�W^����/{zZږu�uX�v�D
��߳绔�������7��Z����7���ڕk(8�� [[?���qpUv��y�_���]���²}!����o���9m`�5[��m��5���(�/~�o����-�y�^�����;�fK�s��.t���瞫R��ۇ�_���TW��yn�L�7M�ұ�l�i����d���կv'k�+�FK�L2�@9�d*Qx-B�ގmM5f�Js��������@�@ �����).�S��uf����ɍ���t���Ä�Fe�0Ĉ���E�A��ʰ��7�t�O2C:���⃉Ԑ�W,;���#�!�����[3�ܮ���{�8�y�##g(~�c� =�����Y����t衽�k����M���1�]|ۙ��:Bǘ��`�}֊��e��iea�30:�P8{q�L�V�껲��+7���g��{��ťIZƙ1�a��@���R/8xwN��Xp�_Z�Z�6>ҋ.ܕο`[Z\�}���gυi߾�n/�+�}�bڿo�m�����$j瞳�X�Yimx���L�+;L���}G�l���x����s�MȏL�䒦��/�s�X����<ώ�fﭥm��2�ٰcV�%w^��s_ ֖��=�3��ڈE�w�z:��rmt8u!�Hq�&�� �m5���`Q������Ε�K�;w���&������G�`���ׇ������w��cǢ�k*����{�=���\��=hb���d��c�K�&8V�wl%؏����w���0mhl���Ǚ��si)�d��k"��57'�Μ���2G;�1k���dSM֎"	�j���s?�s����8_�?��F)��Ϊh
%y�E|_Z��R�-X@M�2g�8��j���h���wZ>�i�Eg\�L���.��0�
fw�u�1��א��pF� ��rSq(>��F��D��]�z�� ,Db�9���w��_��4K2غ\�X�Ԑ�@b�ǉ]G�F,p^ٱ����4X\p���]{�=�ܛ���Ϧ���<|�IO~\��T�ڝBkn/���7�wpݓN0#,���T��|�[���HKۗ�EoOW^uYڱۘ�;kvHM`;]��J���T`|�onM?�����祧=�t��%�\�9Č���QV�D�����Ӿ���}S��������fl�{nK���µ~���� V���i���ih�S7|5�r��5�S��.�e�ԫ�'nӦL"���@�+t0؞�����w��}[/���������v}�=�^�Z��YY�vC��m-���;�}�>����uO�:]xɹn*@��:i?�����:;�*ZZ���7nN��v�k?qՅ�k���pSHi��2��",Uǳ���Nnڿ�7�J7~�oS׮钋/HW_uiZ��w|���&� 4�b���?���a�f�������A��>��?�t�y;�ֽ��y��Y��<T�eS��L�uwJrM'[�d�!b�)l0�}���;  �$e���ou�x�^g��������<զ�m}�(㖡��vk�I@Dx�v��=F�7�҉�[���舜*�Y2���w�c�w�d�r�25p�y�v7C�(���Ka��FdV�YV�����X�DH�Ƭ�A�N>yI���P���*��"�b�����,�}`�1�>ے�*<����=���ƺ�����ϸ:������{�Ys�0@XXr��`���rE9�y(�G>�����t�w�sU��O>+������W�pj�d�f堟��J������o�f���{[��M?0��۞^������Zc���3]J�Rv9��D�Ů}�a��?�����|��I�Ȼ�yOO��S�s�n�Kf�\�R8��������������L�?K�ݷ��ql |iz�~%��ϼ8��Y�z��׺�I�(�L�կ}#������������Q���_���o��0�N��~�f��xT6!][/��[��O�����X&�~�^�^��Wÿ �&�lnM�3�<"���q�������|6����M{|�M�}���[��7�s�s�	%;s7��ܷaZ
� t!撾��/���_ߖ�}��3YL�9'���_�~��ޅö�g�~���X�6[�ϭ�ݟ��~{�䧿��eb�����_}ëҥ�{�=��L��n�� ��l�;�\��/��j�F'?"���l�z�����Nn�U�H�����D!m�������l6�p��}9�-�Z��3p~�*�5Z>���mm�}�<L)�j�i/~�En(?� 3����R�)+�4�a\��&��ᆙA�Y��|�C4�¼�ı�I!�ɟ��������n��
2��Um ܊��9Fu�̈��m�,���ݾ���s�1��N�}������ie��tۭ&�׾��t������jKS;��Fͥ� 	�1����}���M������|���L�_��t���9�r��]��.�[�X�>��/�>�۟Ɗ�b���}0H�x��M|��Ya��	�*nO�z�uS���nL��vȄÂ-�s��>����g~#��k^a,|��q�s��hB=�ή��o�bZ��������a��ᓷ�]g>]���`.9�Ф*ܴ��Z#������_�n�X[pG�n9����䟦�_v�;��3��L@.��u�'>���?�t�@�7X�̯?~���%�=1����gɜ��s�Y93�&ﬤ[~x_z�{?����E깣���t_z��h���ڼo�=A'��,8�h�Z@��u2}�+w��i}������K�Y�??�쬍���������7��`��JkƦo��W�ܟqM-�h�?��Ϥk�{F��1O�}�͝��f���3�:�&,��)�O;A�v^�5��[���o@�=+|��/ RMt��p�?��ϟ1�g	^Q���"ܐ}YF� �F ���O�[��F���َ2L�K+���w=���ȷ���/В�M6��cp3$[���H3=I$�M06�����G?�Q�j 3�;��_�r��}=	�@�H��I�A2VU:�!��Vs�=x�����T�r�	�����z�(zg�mw����~�Ύt�}�|���~�m�o{� x�c�z`-=��aS��H/~ɥ�{\�����c܇:���0=�qW��.�A:��!b����t�}�l��I/�k���.cav��('X�]w�7 YN�\�Tcaw{����ko��>��]隧</]{��y��84��P�m���xMZ?|K"�r��NS�/J���~��������[��_���-=���٦��KLwl����-y�k��ք�!�0پ�"�d�Ԙ�iI��, �k5�}h���K��ړ�x��{�y_|�9i��a�׮����_n >rf� ߷apv�ѭl�[ץ[{w�ZX^��`���M�S�v}z��c���y�����G0ƾ�.{���os{��2]asp�	�U�OI/{�N[{�j݄����Qz�������Y��'<)=��m���*�g":���g���j,���RK���w��Ɩ�t��ķoK�{����9w̕M���m��~� |��!�2f�i�9
ႍ����'?ُ�}^����U8+�Dż���o|cZF��������	����:�`��{�= ��`m���D���iˍ3�'C���R�}�.�8�\�X�*֝7���	��H,J�1�0gl=H���8���JkH4��g�� ˎ�0�hw�)C������8�$r� �
MS�����y�����_�m�/��I�7�*o��u����)�f���$�c�Է{^Z�Ą!y�}gүy�y$l��6�!�xki۲���*=���LO���.��xW(����ܟ|I�'/4�u���.�n0�=���%D����e\�F��^}�3|V�����H{ο��m�1�����Cv���HYIW_�ܴ���;�{�%��/6�Z�ݻ.N�{�����Ҡ;p��ֆ��+�N������v��f��"c�}�����r��@���u����⍴z���򫍑ߞ��w?�g���>���i���t����=+�֧�&d�<P���g�8�oH��zz�ŏI������� ���_~��ߡtnS%�X`>���Dx哯J���-����<-\c������'�N��T^�P�8/p�l�����g��o��w.���g��;�\uͳ��������6pX.�����级>���_�YyT~k������0ը!�0�#��+��}�2(����I�H@�d��s��9��h8�L����a:w��UD��}���������@(F<�D �+;��g=��6���"8
E�5n��g�
&�����d���.��ff�X�Wǅ�������v4sB�l� ԱNv�J̋��^�Nھ��OT�"Z�ӵ�ޖ.X����O	F�I�=�H�];�2}�C�P/K�lm{eg��Q{M������3U߫XFUM���6u�0-�c4,�Jc�;���o�(������ٿ9*킁ނ�gl�ۖWҶ�(���z��⒛P�Fa�E?���"a�Z�<-~y����bJj�d�K��F���a���:��AG�3�����+9�7�ذhs3�cO�q�� �ޘ��E�@t�r���X �Ѹ�����\n;ǎS�5M��������ߎthx��υ�<#*k�vb&|�&��\^X���HR��wβ���!*�fI��{6�6�E�ڗ0u��z���p��g7��j��/,�i��0H����ǀ��	��D0c���i2J���f�q4�'�/�Kc>�7��f�JS�lDՍPsU8GЖ!��髮��q�^B@ ,�p����O|�΂�5!x����c(�3�p�IB�.�c�2�����B�I�P�Vu���#sC�����%7Ex"Bc��#
�5����F�t����sD�{, �� �08�U�v�D�t��*�]�G���މ{��ȹDכ'�g	g�VX��.j2��6q�==��3���Ң����7�j�Q�x�3�6F��p��M���9
Ï��f����
����g7L�+��լ�z�_� �v[��67y�02b>�3#�k�G�NuN
���^���4-�H*�q�l�.�q
/5J�� �g�"�n3'-P��.���Ǿi�e��+@{�5<:��ϻ?O�i4��s!�_\1�p���� >���Z��3�e9���mv���|�x�:������{L{vc��2���Mx�z^��0�%7I!	��� Б�6XH�W�=�sm�p.�^�Jj*�?���I�	oZ�[�#�b�c|��͆$ŐW�m,5b�#���/8�&�S*�G�:Ų��=G�l�_��צ�'D4Ci�¾W���FŨ;���7�JE�}��^��-��0 S���L7�B�Q��6�P&��u2g(��RL^&�'5G��r̓���[�f���L��@Ք�TA�"���ey��\^s��Y=���&��7��sX�d%Ϥ#���d�qΞ�S�F�I��$�.�!y߰�S{!�ը{���+]]��R���L���U��笻^g��j.%9H
��f�E!��Ef�9�?98�zJcAU.��Q����]6��P�zmfϹ�p��� �N��M"Y��P�&��g�7g��q�\gѴ|ϥ�X��x\n���{��)�#B�:O�����:.ܜ$�Ru<>2���g�t-)F>�0��W�x�)��r[�[zd�t�"G1�U�u!��a�؇a��F��D\�Xs<H���`�0f�UL{�uaNf+B�8畣�M�n��N�iʏ��V��*�b��t�wѝM��8�m������K�P҇$#�JI�h�9�!G�	ozϙU�+���:);_:��C���R��%|�k=�^���T��=���uP$�"��!�Cf쀵�NYR����E�i鵅�^��KF&����L�t[��s���n��5*���-s�aS��;]Pns�j���)�$|�^B�r�aO�����'XpG�g5� *z���{�lm��IE�β� � �e:����R2�:ɵu.���z.VD&X��5�&�'�v���GUj�=��hrHk	{<�Wk�i��n^�Qo�4ʢj�q!�M�CNZ��Ir%�f.��I���M��>��p����h �n�
@-׻��0�#{�.4";�N�oI	�x�D�M �֬���1q�""���QvGͽ��l�)����"H.�2�4dL�$��r@�ט�[��0!;���R�o��T����#���2���C3`i")S�i���)��M�t��u״�:����sű�5�Nw��~Y�e"�k��s<qSϠ <+�i&��穩C��y�������۰�:; �IngT�3����=���f]%r�G_c^S�x��47��*�����,CBB��r��=sM.�����(�.��Y�tfdE��6�Ԕ���$�Y�^�jf��M)�
g�.�oM� �� ��2w���E:�Ng<7��2�\���	����!�^
�!^��>�4��dVߝڀg�Xv�G6#��lLcDS�!���Mْ1+f�>1<3D�S��Ĭ������r��*�̖9{M�mU���@���p�Fs��#�jK�n�@�����~�dU����=C�EaX����j��+�h�6��eS7b�����N&7��VPPʑ�C�̒�q�4Rĕ���}�r��\X��ISƱce����*���2�z�9/�6<��Cv�?�l�g��F'��>�s
��$�G6���#�g@S!rŃS��Ռu��V^�`2]�̛�O�z'g���Q�l�.<����KN�0��"C���^��9Fn2��{^�$g��ba*�>q��J�Q�g~�n�/ZC���$W�΍�C�GwT5�N=[*����ts͸)�T:㧤e��k�*MKw֏l fDBv$��~-�[<�2��%���������C;�k�i����`g^�ٍ����p���^������n�*�#�{a�5)LD�� ��0"�̈봰H��<�=/�΂�$�aE���q�e��Ȍԝ��ȩҶ���=Kk
�tHn�$�  ��v�\wOz�o�d�����>Eo���X�d X��r���r�m�y��>F��g�ts��<8IdP���۵�^�-<��	�����٨���B���Y8"ȸ�ŉxo@��Q1�M��XgR��}�����$C���:^"?���gsI؞/{?ޤv��3|�˜�[,�B/���M" �t���\��>��T��Ft����\E��M���~t�ML���7lf�tt�y�8�7�m!u˦��x�S���\5fi.��1�{HGf4�0�]Y	�cz	��n��9���.�Hɶ��7�@PW5�u��,m����VC�y��C�4�����HGd��>��[o�^���ﲍ��,�w��^�|��hG�1P�g2^M��Fڷ�J_��_��ݹ�q��gv�u��-`�ݎW�"��`�5c���ލ�o����`��)wi��<�t[���Kw�������������/~m�T3�k=s֥��͂&r&���<c�;߾՘���!egdٰ�ƖI���r�GUӕ�������r��D�2i &g�i?t���3�MXw�q[��WK����gբ��ah܃W�릛o�݅٨��B�*W�-9h���D7�l��6ގG������ʴ����}�f/���V΀�ٴ��g�
�1�Y(r'�J� ��fW�ą%C��n$�C�	9��7�!{w򵔷�#���i����XA�N,�m$w�͔>�ZβK�o��7�?�#��B���'�Kr��S�1���Q�ěUL��l�
Q򇘵� ��$][m���ǅ���ŏ ����r�ވӀb89�=��m'X��7��8�}��Й���O��~�L�W�{熬�e�z8ruvu�PZ\�xA����� ��>�ZԒ@ƌ�{�e���}���l﷍��[nI��r[�� �9�P�N�A�����%�O}�=�>���h.�C�����Pbp����v[q�{�M\{�A���#/0��b�������?8:��uS@��e1[�5A)OB�;��d��羐r����jb2�%�=�Ո}#E��[�F�~:D��M&W�9S��Yh@���w�|��/ _�2@q}�o6{��>�;���Ye۶�Ё���jj�i�K�n��{䐔�FԬ�X����~��x4I��X�!�N�\k�Z0��=':�):b
��4j"8����S��^��ь��{1�WJ�!67Ɯ1�Gژk��K/;Xxo�D0�^�4VQ�;jZ�$w�岀S�sa�!`�c�SjL=>?���z�hS����rn��x8A�ڜ�&9�id:j%M�a�;H����ZK��VL|�uK[���?�O��G���x�[p7�GM���a�p����Mf��z����7V��q5�~{#��z��Ta��\��0�I!_ل�\���jԉ>��oz��٫aj�7n|�e��a��ٳk�Xp)��3ہ�����/ki�ӧ��X��ςU�@pv����LaD���h�Կ������Y��r���5N=�ǽp����QB�"F�Q�{��*���%�b��5?�X��GS��Gp���'�0��������S鞋w���n��l<R`���Ю�|,�,���@�Ld����n���s���]��Un�w{����Z����XSfԜ{��G��4��(����^���Rs������h�ߏ��9 �@�q* �l��XI�A3��b�0#2�v/��1d��w:!�9�ܖ�N���o���jb�Vj�!� �~�匓ж	=���ϑ�2���8���{G����1�9Nd."��w���8��j�ۼ��s,sq,�u�A�I���h�TY\�@Q8 Sf�F�L����`rصK���6��T���U\x���G�>ua�p1�!J�^�7-ƳՐ���+��x���H�=/��h�?@i3�c1�̘��N���@|+A���JA�vm5�5/a8���hю��=H���1Y9��J���#�K�e*���Y��t�h[f�֖)�ũg�ոWl�
~��s,6�;��a J�8�iB�_�x�hr�iYu��;N�p9����X�D۩�՘r��9��\�����^[�c Ȫ'#�nd�1J�CɄ�* �9r�+�͜S��G�r�a߫�x��	�ˍR�Dݔs/s<�іMц�Ր݇�(%P��TH��yl��؝�8&}��'B�[s�Bu2��p����6��.&+��-bHk�DA\����?"w��[�s�#5��L���#���b{��%_�t���qH��a7V#Ou I@��,�*�VC�+7�\}�Y"� ?��0�}���ĉ>��}��sr2��h]��:����k`���53d���8� �*��QR��:7"u�Ȉ	�Ĕ�b�\O����֖ �+=Uc�
h�#s� .%*/��R�LD^��ƹ)�@P[��XR����%k0a��8�{3q���S\��=q�m�':��$p:��cqXI;;U�hL�s��#��4 F5���0���:�I���d�M���#hSϜN:&����$�P5��Ԙ�����ܔ�Ʃ�	�`�����M��L��27(^s�5^(l�$M��q
 �&P6���ƞ
FTV�TS�8U=����z�k_�R��`��_��t����!�>��O�}�C.T��q*�t�c�j�=����od���Þ<�3?n���xQ"�e/{�W;c��Έ���/y�Ko�7g��Q  �B�/������Ee*�v�, ��(�IsO���/SEÈi�q��#�aI���^L��q�k�����E��7��b�X$�@8&PPY�E?�'=�I��Y���4I<�K�xz�=�)OI��|��ԧ���˿�I���y�s�?���(����ʝg�?��������I�u��W��������I�f����1\MQ|����E^C�أ��1������{ ��C.U�2��DK%lm�0ܡ�XJӛ��*��6��=��t�嗻$�,@�_7�D ����(ō�l���`�0�TJ����C����5,�g�a�L�����O'Oi�qB\ęqf<�" b 2&��U�J?��?�c�d ��i��	�!���gz�`uw��{���2Eo�c�; ��=�y��7���M�Ɯ�p=�6�d�N��Ki�6r�
�4h�y������IP�O~�4I#$��!�)� 3�8^��:8c'�6��1 �4}�+^�7�g~�~�M0pu�PP����A~$�93Ό3����){F��`��׿�����>;;�tXva��x!}��캊C��<���y���M|Qh���&�NEQ����sc��pq�wp�FnRࢸH
�sQ2l���xj-��M�LmF���,���V:k��1; �L2��x�~�����Z�r
%�q];3ΌG�P�����}�5�y�)Z1L�����܄�S?�S���!E:�)8��� ,��"*"Q��`�;ǀ$�XD�:��&d�����jR���b� ���L>mo��I� �0]�$�I���x!9��w�N�����i����X�Vc����[aqL.��n�gƙqf<r��%�e	^��pѾ�����zM]�g��$h��`V��g��2-D;/�rNp �[<�A$C�6���	�I]vJc����;��p�!@G�MIރ�"q���'�C *�	R�/�5;1��b���Yc�A�5����s1�?�3?�Cy@�p�p���g�?�X��1[b����L� ����ڵ�?��\	�k2=/yP��l�;�+0G�#ӄZ����t�UQ�+־�&|ʣ#�bSQ#<��[��x�ށ�2�L�)�q�|N���XP�C�d 1�)�c�m�&��_��_w�x��L�G�>��Ϲq�@��Q���V�*p�錝��83�e�h���a����T �������{y���/Т�  ���A�wԵG�l;H��bBS�#�$��WҴ����pܩ��Y�+:N߉��瞻��7����2R���
n�5���q��7ߗTSz"����;���xA�U�.�G)6�����ԣ�<?���)�i�S7�+UD0w������^o�Xo��\������vѣS�-�H}����K�������F_)X@��W���t�7LqQ�E�ٖE ��M�7'ƫ�f�2�x�F���ٻ�'��EK9�q���1�=N���M������~ћ�E��g���ȉ�Y��thW*��A�}��w)DV�7��Mnfrc�e�Ek��g�ԤF�^�;,��i���k��m~;7y̽��鎿_W['S��c>3N瘷�Ol=�e���"K�c�����.7E��oH/zы�������o�qjj�o� ���
]��H�x�j�����6��P��贿�o
�We�Z��Z.�~�u8��skn=T�Ͽ�)-W\�nP��$V�<C��&A��߀,L��~���CJx
���u�sI��3�ڞ��8��3�f#��4�̩�*��i`��������W�ES�*��)�K#�3��8]c��?�<�Io^�d��u��-N���L�����b��a�Ҷcy�؊(�=��4�A��{D"����r�m���-A�c��锹=w���`��x����=�t1\�b�f�����\��4�T�"1d�����=�d��yX8������Όy8��:����y�{�u[�W��zsQ�<�Pc� l�R4t'):�ku�83ΌS?�懶Y�h�y�8��&<�'��w�=&HH�˷���C/x���2?���W����>�'"	��>�a%��=*��\:S>�U�F�_������M)D�-���\��rp2�K5�Q�1s'���*{EG���������&�8��b�����.[N�Zʠ�j��g�
UΤe�\C��(+��f���j��jG��3�Q��B�c^g�����>�>�6T��?��� F�c�P�� :
��_��+���%��MR��b�ص�+p@X�h%��!�Z��g��oxksĠղ]��<eY�]g�L��AZ_��[5�i�t��p�ܐ��	l�HX.�p�v�vM6c�$��%6�	X�R�e� ~,C�Y��1mne2����g�6oB�wJ�0p��:�������b��c>3N߈���f�Gc�G�����T�:`�����w;�3���%4b0 ����5`�� ��Z��`�2/0�a��e9�%�q8.x�5t�3֝����~ԅ^W�l�U+sm`l0O�}uX��^��Û X_Ib�
��
�}�P$1w�,��!;���m�]~�b�T�GP-�m��)��+J�#�i#cq��"K�c����ek
�9�Òs7\�Mg��,���3��3�4��bs�&z4s��z@�}1ѱu*2WE�0;���o87��%��5@�$0�2X~���*���1Ҧ{�]������5d�I�i�\vG��	
�$1��(���?HW����(�zh�n*'^ �j����3��"@��"�H��*!S7H�5�Zbk@� l*+���/v�ü<�R%�;�1uʀ	* �1l&a�*���
o/�tS�-���t3�ٙ��1m�әqf��!�Nb�G�cq�EU^�SU>��p���'{���wyf�.˱j�@Kam�0��`�I�>Eq� ��5���\��s�po��焩�Qi	�rFk`C���|��_N?��t��d�ét��3��S 5�����_���}2e_Aa��+8�G>��h�X 7�:��ɐab��'��>�չ��&[f�t8�,�ic�PZ^��h������x#M0����,E�Y�1����pL��N�tf=��������P�6������S9A��=����L���L�G֦��0�ΜxM��暡g��Bճ[���u*���%�ߏ�i9�֔3&��S�RϺ(6T�QlI����[�T����Q���\߉eY�7y���b�����o�yf�V�<[�}F߈�I���h>�-.��0�;Q]��6�G��BW�����ǵ4o}i�D���*���x���Ҍ��Km�M���	u�͂1� �	+�-�װMS2�h�M�>���2u�NVۛd�`����>������!҉UGX7�E�bPzng���~��n<���zP*���u&���"Rڳ��c�����`�t�[V�k���0{�ũ�����d���R��U����Pw=�Mҳ���	���`9��Ua�f�<|(�y��k4W��m�3��D��6��ɟSP3��kk.cXN;����q��0DE��,"���Q��q�ц(A�s��qbcƨZ�dc�dLT�E0�wb�,�������lϟ%�d��rZ�
i����k$�g?����磹��IQ����9"��ׁ����j�;�u��p���k�5'���	J� S�G���I怈����b06���ߔH�%0)��������	�;h�C��N�8j�e�=U9�����v�^z�S�꓃���r�jE�`q21 0��=��J�j)�Z�)<�X0�I��j������l�?h$�(��I����sv�z����0���4Y7 6��v�^Y��tO�p�KȞ��~z��Ҏ�.rޘ��λ�I��E1sv(�$n�MϠ%��_�U�aH����<��z��Њ��^��o�TF[[Խ�Z�uEO��'Q�n3�M�v[=k�|E�C�MM܌�P�5��ⳬS�[���j�<T�J�V��GdB����D ��� MZQC�@=G�T��U�a�1�I�K�����c$�T�ڶ����h�k�<\l�B>J�ҵpm@59�t�|����<��`Eh@U
S�	������o��?7�#!%�*�V:�q�*j�lc�䅼h�nf�D(�ݻ�A�e)y�Z`L��j ��&H\n��b�I=5ew2e�d��L����������mS�a:�3\�����0m�Hc�i�L�o�;�L��1?$n����z]S��:�ԫ�>�*�Yl��`p=<lm渨�����.��{b~����o/J�#1a͹j��D�>��f��jck��Y�X�|Qx�"Lb�z�\" k=H��њP�n	3�(x,�{�f���	7�Pe�X�@�)Е��c��L	F��ya��9��F�>/� �}VM4|F�s]7�M;ZC�5�sH�E!x2� [�Yb�c߸H�tj��� �-�^aN�_�������7��y�w�|E�TSq��xtsD�)�d�OV��^���Ƃ*�M�t��܄<7s0^-ˈ�$Q�e0	T�GRi��q�yO���g4.�gK��b4d��c2flG6�P0 .�1f�I��ii��a|Ua��h@�En���Y/���{�nV^�s��$�z���,7f������ʓ��`>����N�P��h��L `��uIeBj��GtrD6�g��1�R#�H�&�X5jM�髽�/�f��\Q;�J�om.]s�=��hֶ�1�:�3����Q����ɼ!����(��֠��.^׫=5�v�A\x"㎎>�qt �[_�2��������K�A�F��/ӵ�=�t :�	�C#�<�u�s��^�k��jFDavl�i�>�z�2ؕȎ�v3��Q7��Ҡ���=(?�
*��D��ő��a��E�h3YZ�L���5ǖ=O\�Q��h#/��*��Be�W�lA�vX�^����~�<�*���ʩ�%��Pc-��0e�,<dc��R[���b޸g1Xݣ�����Rs��m����ܺOƑؖ����D{�
�G0��#��Jz֑-���)@����5�_	(��~�di[0�L#�D�b�1����������"���~#co3F���Z,�=�q^%����H�p$տ�^۔��q�g�&2Ui���ccp�cQ9Q�eQ��פg�\D|���N W@�-�����x��=#	�h�kk���p��V��B7,<�A����ͤ?L�����T�B):,Z���iqkB��8��c�6H���&XFcy9gj�_~�1��������
�#T��Sy���T�̀Aẜ4N��ɣ& ��Ttlsv���y�����]6�v�T/چ���0�5�V���5�,@�T��E+�)՜��(�E��&&�+۶Y4*m��Y��)���H�"�^ڂ�k�����F�?F�(
�m�՚��x���<en�YM�X�����^P	 1j�p�f���5q�<j\�b��]ku=Q(�AYj{M귀���6ؗ1��D�� k�k�ه��_p��ڋ���Ks�&��7�)��s��k���#�(��υ=*&K��f��ؽ��Ә@;lʙ�%�WLL�Ɇ���ʪ���V�d��MK����~�Y2����<�ԫ|;e��~�I �669���ML0�k�m \t��r��oRx�v~�H�$J���.a�ndw�m����[�M���juu�Ȝ��	���?7=���{|��Ճ�7�;���cr^g_��������~&��{ -�=%c2��l��;�W�������=�g"n�8X�lr���[F�%������g?�m�b�Qk��]���Cj��72�ig�V%�Mt�I�s<� q�j�6B��vZ�A�^���CmU��(��@0���2ma�� ��ԧ|>�k��>6!ҷ�76�z�����tŕO�s��.�����'n�tZ�=�|b� 	��]=��\͢\d���(������F�C��랢�"ڡ�}��s\=��@����A�	��)tO�c��?�HĮ8�G[3�aװ �ș�b6k!4�����4��u��ۖ����I������P��a�9�f���΄�Xۢȅv�����\����l��.80�;������NDWTv9��1ݾ���$8��a��G}5�cM܎'n�÷[�O�:A�c�#ۈk�i�9{Үm;�D޾���Y��i8)����7��ඥt�TK��L�F��P��?�d;��h5�}�Y�
WRJ��mz���"� O�Es�g)W}c���L/����F5��c#��~��
9��%��h�I��1�F�$��E���(� ��Ħ�&�/ ����v��J`�	׳��3�]�3'%�������{}c--��H;�9�C&K"q��c��ʆ��8d�dt�������	���}��~>Cy[�k.�i�N���=�ԥ=�~�N-�����5F�������8M5}Đh�o�i��{m�,~�mW�Y2~&���L<'2�nY�ug�Ņ�-�������w��BtDck�EWgV�����N���q��#n�u$����M�	�i�$8֘�0`g�|	'�Ԧ�T#�dݴ<�s&�D�ƺo�����IAH�r7�5�5�6�B�Ū݇��n�>V���bw�����L���Hy]���T#��V"V�!}V&(9��I�#�p���}@�]�Ҫ��F�/;v:�� SL����C�E�C�I��X}&F=�L�:Eژ��ӛ���+�w�kB���Ę2�Au�ر�E\;8F6*| <�:'v*�j���
5�l�4�ߢ���#"���8>/=1���F�����8���'q���V?z��a�K���6n�ܱ-Б-�5c�K�m����ma��1������6����պo��b�|/D���ӛ�dUiۤ�����*6�1�8���Y�x�+��U�y�LK�rw���{{Z@�3���k�bv���7ꑳ�����%cT�9�Y�Q8V�AZ��1����<�����z���.b1Z��K�f�A�ًRP����� �z:F����,#������D�Y@ -u[ -�G�G��f��0&	�s�Ĥ)�����N~��][���!�nH0a:H��0�~h��|���&�T-6�1p�%�r������N�+����T��ZN���%��69�"����qޣ3.fk�7���':�i�� �g��9r�y�}�d��|�ќ?�D�#yH%��$��g,uyq�H0�2���Tum�ox,������=.�66UՊ΂�������0S ;�vw�V�c�À�t�}nBź�)�~(���zm�~�ϧÇ�i>���n�X��?�=�DK��=����D�`����n�O���O�s�O��S�� ��qd�n�8娐�]aal6JR�C����8�8.��WLWj����qS<qt.iHȡ%{���� 5������j(�����)�#��R��_w5i@�l�W^'���L޽�,��se��;�Pdi����l�84J��ݟ�n�u���߀�Wd��J���&�����aƵ��IZ�,����lJ��M�8��h���*��ˁm��j�J�m������T�~�wƹzjL� ��v��0}�;?Hw--xDDQ�p���jºJR	�m�.���V��`ˁ1սE�ƌʅ����!��� P��Z�W�M|�}}uZ��ҶA?�����;�L�{J��ô`l��R��ᎪQZ��9�7�\YN��]��z�Kd�7��q�s���n���-A�����t���0!1FEN��V��bYb�����̥���f|�8�,%��?�߀	M_N'S�;��~�@�L���p1@���y1��1�k�u�E֗��7�2���ם���\7L�*�;4�nB{����u���0�� ����`j�"'��lmM���v7���:5����nn��A<2X���p���)2�4'��ؠ�bw�O�7��"���Nt|O�����y���cl	���W'ɀ�$UN�}�xg�{,�I����e{؛����e[#��5�T/o�i���~���mE �nM�0��RNY.l3q�ޟj`�ks6��U�R�D��y����ɚ������;��=Ʋ���� X�f�kc��&����s�6��)��Z��_�q洸�O��Y��tNZ�C�QvTm>1���L4��]�,�c!1W�d����G �8��4�}�h#Î��y�M��L�Tbև°\(%�O9O�f(?W�U	&�$0������y2���a�V�[���iLd�{���y"�a��>����l>��Qu�rB�k)fi�1r��]��m����_��1Z���d맿[�-�o�	��G��9���6o���u��9��u���Qi��6�:�%�p���X��X	��G��l�:)���56��iNm̅�aSpP��&Y�����W��:�me�iTO�O���Dc`�s&��4ZM]��^�M8��,����#���B�Ŕ�U�����h���+;R����b�	�S<����S,*߶�	�b2Cj|���"C�"@�衎!Q����~R���c�� Gl;�,#�ơ�-%X̛��� u�a���A�P≢�Wl�1m��Fk8�kꘖR�h�l�u?��Ꙫ��0���$�'o����sM�T�"�3/K�w-��&�l��Hc��N�<dGG��(���4�c�fz}�#�DƑ�b4{Ź�@|*�tsD��^0�����D�m���U<�ei���:�N7~jT��&�v�l��V�G@d�!v7���V��no�`���մ9h�#�Rj��:+���x��r�������L�u�����H�_��fd��c�w��:����9�W�"��F��v����x���!�X	,���G��s�Q��\����$�(,�������	��E#^[,����y�n�+���{�N�q���	]н0Ѧ���'@����5@�K���Ԍ�򣻝�y6��Ud'���L�4�_�I�6�T�H�GS��ޓ��dAj����Ɍy ���^Lw�Sk�E��u���(-���PG_\�c@5N�y��T�"!�^�R��{9P\27�� �%���Oa@��dRT�T��Yu�Qy|-5T����^/�ncuc����:�~ʙd�T9!y��o 	��M�J��P�G�p�I��י����kg��l;6Y�Y�hc�� 7jc6�@b��N��"��=�(���,3II�:!a�d�6L�Ʃ�6]1�*͗�S@!0�RI	�lJa�C��6#��x���ڶ�vWLmg�"/2(*�`�fo�λ.]s.�+1�NS�I6��	���2,I�1�h?h/�Fɸ���z�a53KW�
w��S ڪ��w6��Dj��Cg�$�ǹ�(N�ͯ↹�X��H ȏb��~�����v��u]J��?�*mb�*&{t��^�$p�VY�`��Z�D�����b������<1��%&��6h�+��v�?-x�*�$�� $��U�G6&�������ƍէbH���3�4?LJ,����nm��q#����z�<���
�����&B"'��D��F-7H��\e
���2[�,4����&��M�I���d�8R������h��_m�ڦ���^6,˄@�͗,�n'�D�*�=��k�����{�`�f�I����7Y�o3�x�v�!&s|G
S��<���B,�?��3d��gu�z�h#�_���:�NZ�׹w���JA@W�����>K�M�%��
LU�ak#[� .����� ��w&^d���=:n#~8FDD�SL�j�蠋�(͙b�e_>��5���I [6��p,��H�3l�d`r="s�Y*dN L�4��Q5�P� �؄��I�	��� ��-�6L:�L�w|'���7\�"N��p4L+���F���~�9'@��.ʄ�D1e�@�M�K��X4nr-T�`_�җza ���}��.�X\1uV���e��JX����[4	ިsҘt<>���Ÿ��Q�:�d
�\ �.TfpV�g�b�d4���"�o��!���Wm�x�0Pi�k�Gg��c�7�=\{z�ؘ��y�s�u���=�s/< �c����a�3�换�:HsUx	?%^H�V�39͢SL�}�*Tx��N��<����Jh��s����ў}$[�Q�E��A����V�v�C!:y�J�W(B!���Nm@a��%���4�Rf�n�*�Z)��i4��J��:9i���������q�ur4=;�A,+���B̈�&#���ﴝ[�ʄe��is��U�?�J�߰c�븬IՕQE?��MI�`*�I �P��1D��K/ubI�a�tyw��D��l�3��n�U���$g��];��Wz�>҃I��Z찡,)����{ 'L��Efx��� .��2/MX�z�!�uW�ut8Z�{Ǟ����]w���;��{�ңO�(T�~;�,�n�u�����Jc��Ļ9���F�cˈŗ2�N�5OS&��6�2��#�i�c�� <�@���vO&��?��k�d���Yp��}əyUO�j�I��[͊��ȅy��h�P���Z��<g͑���y�g�bF���h�����o����J�D/��H)�C��h���Ѱ�.l�wsrVd�J�&�nl��=ת��Z�s�x�Ɠ��̩����9/SN��Uk"th{�u`*�L�2���O�y���[a͋��U�pL̐����Dm�\1��_��w�t���������Z_҆b�r��A�=+��Z�� ^1t�h�`@͹�.�@ c�f�TS�r�0�tSD��9>�E>���M�|�3��=P_m�5Z�|I��7`̀0�O�yL1)�T�0��"���?�gΆaҔ���=��H=y��$i��E����4�>9��(��=lz�!��*wZ��o�!��p=3٢�馆9:[�x�*兺�i�ôL�1��U5%�yO宭~a�gp��r1�ln�Vؽa��k���4*5�M6�Ϯ#^��mA-nsU������_��X ������<�)Ô]8�T#@�TN�p1�-�-^S}	=�y#:��(�I��n��U$f�Ţ3�OF4U�m����ǐ�-�*�2w4n
[���A���u��l�{v$x����Mc������8�Ԧ(%R�b�k�-ΐ�F���A>��Κ���[�>'��aqi0��5�}�vHEgf4G��(��C�x�|T�b�v����e���$�b��4� �8h֊?���PR�PÆa�M�UeF�b�0:α5�t��b���Ƕ���~���'x㼃��E�쓣�ǐ4�i����dw�_��88�q��ȯMHf�O��O��O{K$���o}�mx&�caC>�M��lBm��ZJÜ=t�9��A��p}H)�4 �L���Z��rvR�+��xQϣ&(�C���c4��{�v���fZ����V�@?,�P6�ҍq���߇+[���C�l�~.�B��}u��3���������>�q��w ٰ��qb�E�K��\�8T�W�P�{bќ�؊�@o+O�l�1ck�sN��b�v14��u v�k�|���Mm �JP����t�N�mJ�FR2�χ�r��gK�� ����p�M�����][O%�b>�u_�y��.��i�y��z�F_4)�N*&����8}�C�|h��ƽ�&4X%��)�1��Nt�� b4�|��^�����p�~t\WK#=?٤�7&X0X��7qM�u�>��P��z���1Os��ԛ#tA�ⰝB͑(\<,��y�*Oi�Ǎ�k�j`�H!l��^{�Ԇ, M2��t�M�]�~x�9������l;}�:JٹAhW�υػ�4�:����g>5��{G�G�Ɣ���{�d�pZ�i���M@�Q{Y�\�,|�(h�-��>s�b`@oB��!7�`�@-�i��ձ�w��;M�[�2�����0}�4�Ʈ��Թ��&�'`�)�h�ąцmdJ�7�i�;�e�.�5=�6�!j��LE��:�1BE�]�o/�dX<�;�V�X��~���u-mm��[�&p�K폩�*D�cE�m��+�q����?��7��j���E�:��8�4�ά��-�e�6F�`~�F��ɨ㭳&�OxM�Í�!��J�]T�L}e'������\rI��)4�̚��[Qsh�6�����g�"Lt�A�mW�;���zo��]s��*�$����7�ɳQv&Z4ׇ)��DS���ֱ�U)�s�q�O%���\7?u}�R�� <��~2�Z���:�m�V�7~��n�X0�{eI��#�M�D %)�lXn
�D-X&]]
����w�ˁV=Q#x0������XY�9��`?���A�Bw2ؠz\|�%�=g�Vb`���8�(�R�6�Z�,�(|�0?�[��f���+uw��g_l����R���{�t]=����h���͹�ۻq��c9u�=?-����Ѐ����f�O�A�T6��}C��{��k!=ɀڱ֣*RZڶ-]x��q�\<5GD�AJ���j�ʆ�EK�L,p��DV�A,3o��*'�5�x���4�bW}Ւ����2���lLE���)�)�9�Z[јp:M�a^����0�8x8��ƺn�ޝvM��R�J��봲dp��!���j��!�y�!��`�~O|�h9USv�����bP�<7��s[�;}/o߾��J��P��CM �φ=�e���w<CRp���ɚ� �u�z�f�Bz<D: ���������V�4�V��4�;�U�
J�z.:c7v��b+u����\�zt���+��Jm@= �/�ls���NX�ֆgp\�6R�̓��IT,#���>,���<�y@[�^�p��|�/-m706)l��ǾKҒTɲv@��L�(;�_�C<�t[&�!5aOEV7�\%�fٔ�d3Un��̮I��,L��t�������Ҏ��Vnj ���������Â�ۢ<�p�2F�X�=����x�׆�g_�3�k�N[-�_Ӊ/�_a��h<��zի������b��y	��M����Ǝ���Ƹ���Pg-q<�1�VD��Ą�cFN�R���ņqİ�c#�����H@�{�1���Z��G>��gs}#�B�S���0��t�B����4�)��ͼ�YX`���d��VǦA��)�dߙ�����wsY�����&��h�Mh�^g*���2�u��D��J��##b4J�d���W�WݎKQ|��F�_��z/��)Z6m������1fz�&�+�w;R���=�*�T���(�6����i �Q�����������t"7�»g�]�*[1�JЈ�|���&��;y��E�Z4f����/��/��U�w��Ƅ�������Ռ��,:�x��Ԅ����,7�gΑt���"�D�v�q�^�d�n"�5^��].�=u�Q�%z�SVY�,M&j^�E� ]4@g�k��t���Rw����NZ$��>O�:�l#;����a��`�k%{��D����dV�K�7�ܤeD#�Q�����%&u;Y!F>�ϭ��ܡ�c$�W��@�k�@�=8f��d���	��O#�@��Z��f�H��/��<�ǔ�̟}so�L��\J��d�x�4�Uڜ�:�����»/ w����S�{� �N�O�7\�%��漺c	ӹ��8��8����@�<�W����^���?�A�|���p
 g)�J �u��i�J�H��	��c��M�O�9"�BMg1��`��6��K</�=n�Ȣ�jL,�E����t^}��n7��G?�̤��o�V��?�c�H&Z^q��F�͖6=���m(*�Ԩx9�l����u9�B�<C�3����^쎿�|�QAP|��i����g����,?t���qӪi�X�r��QZ�.�=,�Н��۲�86�3�̞�&4������o9K�Öp�=*\P�|�|%�E:̋z���Q���'A�.�.��-��R��[�/�4�yf�h���%tt_ڴ�L�:�K�����I�'w8I�X�g7�����L�Ns�\�C�x�.,j~ǃړ��o�Zݸ���x��,}��ż +��a�~����{i�<G�V�g�o���-F��GX���7�A�LII�-;'t�Gi�9�	kZq�ZZ,9 ��Yeɟ���1�ͅS�6Bm\&P^c��̚�����o~�g�D'���
��^���ڧ,A�h�K]z��=�n�s�$%�Λ(;U&I��p��w�kE�Ջ��zS��'^���v!��n���t�Ъ�g��Toq�$�&�y��=���-��>��1Eԓ���H���~�k���yc��s��`S���v��
��9ڀ�F�^�"�g9/�}���ϫ�ql
ӈ�&��)}?ޫ�RM;?�Fvg�����L$��g�M�lM�����{W���4(�Q�m���A�Q&lQi���%��}ዼ�e� �o�,�ʠ"����4qq��1&Ј!�Mws����C��uߟ]ߺήڻ�34���tU�}���~��o�L�͂�e���%�}w�Y�l���#�_�ş�m=?� ����;�JzH:nS^�G��f��m���꺧e��X@��>T�	��I}j=��'�i�K� F�*�[K�1.�H�"`�#�=�;-��Ս�S� �7/��J9�tL�]�=���:���j��h���§�?��W}�W����� �l���=Z�a-�*b�����P��А�I9o�sp�3$C���%v�9
6j���YHK�cx�+W�){�=��ǚw���}�io�:d��VN1a�ӈ?����5f1-J� ��u}�����8�1�ڎ\�1tP�k���ph�f���h߻`r< ����1����ZF�����@�7�ɧ���y��9�G�gl-{+4q��x�w���K�?�5l#)	��d���7�Q_����m~�����?�áF� �����-�j�Z�	�3��w�l
�E1�Fx~�NjEc*�S-�������,�������(�n�A�,�n�<�ƪC������,�^���?��r�1�1�a���@��k0�<c<�}A0�LdDk"c��D�0��5�yM�,Lt�-��|�:9��ps���
/ԍ{���%�s\ �L���߫s1�k�ZM��v�=���:4�|��=~m�	>�ȣ}Vނ��*am�o�$(����� ]��DR@ee�עд��L���M��s->��S��a�Vh߸�bΥ�+�@�i�V�㈾w��L&�X��|&�'�-:����8z�� k�ױ��(���h�=Jm�[�='������c��1]ڥ�}%������������gǏ�e���0�X�H��������{��җ�z׻�W��U��^����BQ��:��g:o���q�d$�ϩf�!��x.��|��h<����Ɂ�s� �O&7�a�j���y��"i�9}�>�:4a&:x��v�=��=%���:xC��?���q�1ji��'e<�$��j���>��p��Ӳ�r;l�9��F�h?�X�z��Ds�-?WP���1Y��QےSЄ�x�䕽�g���|ڧ/O�>;oww�L�@Ts��#uw<�Q8�_�K�z�C���!L���.��km���\�7kx$Ր���i���uԴV�D25�!�$�M(��Arۚ�j��&9�右ԧ��&��Y=����ܝ%�G�8Q4Kj��К�h�Mb	UcK���I��Ej�q���ӂ�j�7^?S���}
D� �l�%�@t�l��؏�N;���4��x��;�A��a�CA
l:�Zt 7@ȿ����1�wc���xy��έ�,+?QeNy:W�T��A����tB~��4#t��9�����P L:~��++�k�d��%l��󶯐F=��bҁl7q;�q�N��ϊ�eT��+�Ep��{�찱h{��h(�Px{�U��bqXwb~Ѓ<�=�Bq��;��Z��p�l�V��ս�����xf�+����o�����u2�E�䲬e򢂗א����w�m�L��woHmE���JE$�;񼎜5���j��<���g֒�s���¡W^��J��h�v�ԕ�;�I*�}��M�����1�<w69���4ۏ����;/}�{1�q�!�`�h/�%�W��v��3t��*<�5nҿ`�t�%T	 0A,���J��i��dMx��Tc;+� �^F�X|�+^Z �����b��H��9��z�iDB=hh�uZ�	!��M�T8a7_t���/���MozS�����z����LQ��jٞ�w^=婟��M�>O~��.���uZ�b�M�	�ޏ�&͕�I�����.�&<޽��~0j�ߠ@_�}���{�Gy��j�m8]�:���e �յ� �~}/�����ﷇ%���b*�e*m��LV�{�}�V�Ϭe�����;�ɽ�N����'}��<n������9�M�-"���֠u/4�3�o����MGM}LD�g�g���~پe�|���򓰧r���w�^	��G.<�>f��$�>j�_��=Kz/�˒����0w�F }��8yv��P�x���ȏ�HyBW��ۿ�` �,kS���Ll8�+�`]�h�j����x�Mr��K1}����i�l��F�0Ԉ��-@�p�7m>��Z��08՜h :�����9�A�\(4��_X.╯|e�v��_����Mf��|�ה8a�w�աL�t�!�Xj�P���o/IT�"�c���"���m����H����E��P���nF��{:��4�+�t��Wڍ{Q�`^���)4���1ͥ���̛e�qn��/[��2Z�N�^��j_d/~��/9m�� HH�0�8��YZ��I�i�b�2��h!3�.�k���~˷|KI�b�������_����q���Z�8H0#����#iK5^1�s��(�;ڊks'�:���S1h/<:�4��0�c6�/� �0�y_�З �f��	W���X���r�(/��hDk ���[�Z8 �6�5X�h ��6���P4�-����/�i�&&G8/N%TƗ6���(lo�y��h;�Q��+���ލY��P�	J�ٞ;�5�5����.٨�[����KS��C�:�/��m~����e;�Ns�C�oM#��VǶ��9�~��eJM�b;-@���D�Mjg���?�Lk��U����#:ɚ�ʦt�?������</Z1|1QS�IF�Xl�yL�.�n�������n�c���h���~���Hџ�n'eXSDK��~o�-��xz�9�yn����U@5�Qn�tP�����AepM�BY�$�O�tb%b�"&��m(�#@�Fռ���a֧E\�(�X�Nh�=G�$��L�}�Jj�Bo�8�+�X�o/i�MS2�F@_�z_�1&K��q��@g5,%��k��6j���tr&��[ṿ��9���~n�:�l���f���f��c���|�*R�s���T�N��:�Rt�3��"qȓ���F�3?�3P���"w�A��:d���2��5f�N��҅k��v"<ҡ�mw��s�E���������~��>�O%��s��9�QXa0G [�4n�B^����ĺA��q6�f�GkF[��a��m���Ȟ�zm���J�-��1��b����%;���(�4����h�.�6�������<���L����G�5ړ&�0Q۾OF��IC�)��t�3�U[�di� �����'�(J���SN��c\>�
Se�c3U=��{�iE��v)/���X�k��et�d�&< #��%��ǝI������'A��zqqʸ��X|뫨����v����%�΃a
�����8P��z��Zx`V!~Ҙ��h��2��f<� �f�3L��c���Vɧ���������a:��߸D?L�^�-�/��{p�H�f<�U���z�Rf���Jv�25rѧ1�b'[)������Ak�{�5C�E/�C�r���]0�H)�v Ϊ���d6��A�+�*C���=L����0�Z6Q��M��K��,������OxN�b@�H�YZ��BQ���8���F�P�_��Хh�p��x$Z�֋�#JC���fm���a��br��,$�y(��)��B�~���8��|�s�j���%����3�+�n���9�`8�㏼[֝��u��M�މ
)��P����Ė�:g}�>�3���[�Þq�E30l pI�q�ŰS�
����WO϶��%p�=]X�e���	_�����r+���Y#�qյ������I**���T��SW[q�G�s�	̂ߑ���6�Ęm~�������6܏W��CJ��35�<��qԁY`ֹ�9m`Gٔo���C�?�UN����S�=�Gn�r�͵�5�>�f���2n@$�U�m�����0����
���Y�*��*H��Kj���gL�I���Jl!�����"��+�q��Җl4����Í�q6lٛ��sQ6U,!-�i�ϕKI�a)�c�5��4SգNЧ�r���;��>{Ϻ�p��!eF=���xnk�x�*ǷU��T��y�kA����P\�7>��ris�NI�	E�@;�O���	 ��9��g֥���!:��5�����3�#�d�C�ס�}`�:�Ǉ�qR+u�T���d�)rKj�5a.@g���l��$鷋�,'ʃ�ڎx����)1F?��	���5{V"ߢY2��t�O;-{�!fK(��]a�rl��#�mn�܉�o�yE����cW�����)��sM',�4ڥr��γ�x�JTt�o�(��Ӷ=ǳH�Ů�N^��]^:��c�T��������q��,0�K�?��w̝Sr�����>I��G�N<��?h�y+��ޠ�V�w+�![�崒���~�ߗ-���4��΢m6�|: �z�W�M+<����V����!u�S�~����I
�I�$��5g�4��ٖ���rF	̫�n���~�����RGc(�FU��~��wV�
M�,@|r����b#�$ d~.�m�(���滕�|��y�vS��*�=��׶�x�ss���5�+	���^u����oAz+[yb�y��e�����d�9�xf^8#�ڱ�f�me+[�����8+�x֬R7Q/R��i7�};�3k�.�q���)�-'���<qe�OhU�^�y���*���	�N���n)H1ۛ���>{��|�Q!q�f�el^Vg2hN��5Ӕ���6_�Xd�#��B��4P���m�t[9��s|���*ӯ�`�
�O9)�,���DZ�s���\r��N�:���C$�`��kȝFΛ�h�� �i��I0�9��w�sS�3� 3��td��c�M�����='\J<��O��Mg����+[���zG1���������9��[X�
jf�X@�x�6�ŧ�\�L��CLY��j9S\�	�)'i%�����}c�yN�e�b{�k�Tw��϶V�v�=�ռ2=xUM�z�;	\3�vG#Y��y���!�o��3=9ے���Z�s/::��r����ֿ1}��`�G��Ӿ�uuz�v�;Z�԰�O�[Y�F��Ew�����+��Ȁ��C�bn��dCԓ��6<�n���f�]F_�
���� |�y�8�:���R�:�cV�����LA��%�]�o�9ۮ��vzזF��*P>�O�`O3vΫIg�Zֵ3����cb�J ���Z�f蚒L:��ӁUVU�������pV���R�٨�����bSv�����G�8_W��Q`��Ǽ8`�N�!_���`�bd�d�[�˕�MZ��t�ֳ��|�C*�������x��ǣ�2)kJ�,�L9	���]{�8�D�ʸr��IB�����.I�X��8z'���ˤiR����u�[��B��Y��ZH���w05]��������(u#����N�v
��W�."�[*3ۚ����|:m�����H���~g�8ǻe��g?��e�^��GTw&
�%.)�p��=��x�41�G�����5A�/��//�Q9�FB԰���J/�&���i��d�{M7�,̀��Ȫ���4A}N~2���� �-s�%�U�A`�
��֝+�iL�֌�ɂBtn�$����Os�ӊ��|/bXn>�q�VV������g�
l�6�#���T��d&xC�]�Q��1�����e8�vvڡ:P�}4�\L�|v���^���y����BV%�C�MHV6��8jx��g�8��]3���W}U���5��k_�ڢU��~o���		`#TB�o�x�UZh=iO#5�X�l^7�s���6Wq��-w��=��K��w�d?���bCaj�J��~�p.B�c�t�*Mv��c>�Rp�0U�jk�*��Ɗ��������+|��e��?��?-@��(s�-Q��������F��=�tI�mt� ��؎x6���lY������K��-���4��<�J���'�̆}��^_Zg���AL�p}@͘	)���v�s<��NnX����ҳR�9�4�yMM��4�$�z^:��kgIĴ�r���E0�m2��ww�I�Y�d����}�Y7�Wi�g�\��������h��'4�t�%��ri�_6��P��$:��������= �`}s}�oJ��:}Ԧi.A��Jw�	�N�CǰR����̧����R�݊���N�Gx94TL^��/yg7
u ������-��_�x�7U�9���lYM#
�4$�cʥu���x��G�e�H~�����owQ�3��e��ŹG���zCG�Pw����7�U���w����y�i�o�9_;p�x�\���_�=��X��F�<Q����;w���j�75Ԛ�Y5�7q��ǿ�����:Kd�Eܟ��`Q� N4Y6����_��%�HG����Х/y�K��P����(vL>�x�q�A��<�X�+��+E�ĺ�6�:B)��s�^��3>�h�t�������_~xٱ5#��/�Ơ4 Z1+��ԅQ���c?�cE�������5�{<q,�����tXzVW˨�ض~���ge�N6�/v�M7GlY��Lg��рp���-F]�-��>�V�)\^S�zQ6���iL���x���	��l�Xn�Yvʘ \��&`s�L�Fv�6�^�ٕ��b���^�κw=�w��)�=Yx�S��;C��E
�!���G������@�����.)8:X\��?s˘�l�c��������n�)~�J.()�$�%�[K_���
YJV%��5��?�3N_��]m�F��>�s��������׽��2�%�k�7ύs�x�[�R��s"`;%���/,�g�b ���MHݐ�cxfϷP<�>�_��]��3�\��~Y��\h/l��áŲ
 �L4M*�&C9�2��5�8��b�¯Q�cJ�-G�dr}���+t�7}�7�p�n� ��|���>�w��Ґ��W���/;-�^5;��y7��zf���x/'��k�:��4�vV��Ѽ�9[܏5�3-G�_]�X���w�����~��q�i�������4%���]:&�Bq��N��?[.<�fm�N���:ۦ��6�� yw^0i�]m������,���e���a�q������������rZ: )!��DY�?���B�o��ļ���6E����j�*HI
RF%����J:�yf3}���v'�|n2̎���:Z���Ԏ�Fay=#r�C��ъѦ�+�jX���.8N��\�F���<��4�м���备?��惥G�4�<
/�>N��4.Z1�n��G�����ſ�e C�9\�E�x��ye�i�@��݃י���ʻ;�d0�H�{������®C
p��8��i�N#�ǃ���Ԇ���>���]���+�9$â�@��]>��� �N[���f��כ��N���V�!C����u�$w8N� Iڒ����zf,��Ay5n5����C���h�Z��|9�w�n��N���]��M~ү�- @�~B����]m��=5������:��J8�981g9�t�����__@���/��|M�������=yN�%�{��9p���X&�:F3��4�
$44(N:�o�UЇ�@�pV�*؁�����}ۣ�f��~gRUx���ܣ*�s�Hh��X=��̎1\�kp]V#���X�8����1���t��_G��L�N�m��k
p�A�l� �u���ɴy���Y����On��>�\��)��J:�n4���f�j7h�,�\2ل�/FJۃ��M���#�8��a��Y�ni�䈻����W��z������>�i��d�e���Q;�l�KS���a�8q���1��d2��kq}���o~s1ɐ�]l�@r�����jS9/X��"�����T�k5U�Ѽ��C&@e�WF� �=�P���8)#��r���� ����/��������.�>	@73��*����:�ZY����H�r/>�	^l����k�q~�tD{p�i��Og�x0CC�/������;�Q��2H���n�t�����1��A�P��4���e8��t�<�q�7���{�o���sԻ��2{��g~O����o?e�\ߟ�ĕѸ{����f|�����|�k˅����\�
�:�����y8f6�μt굝	����{�m���zj��]��|b7Jz���μ���Kʹ�׉Tm�֜焳�4����O�����51�c�#�a0�%���ó�w�$}PG�lz�����ڣs�߇
�o�D5��\t�Ч(C��I"R�ab���y<������*��+^�l�5쳨ȩ4�ǻ�#r^h�!�ͻo���B�uhC���]��`ؓ������9�;�Q�K���R3���0$)�U5	����1܄I���te��il&4�<&/��{L��FE�̣%��	Z`�v���9�yN�_���=�����z3z�Ϛ��?Ҍ��E���pʝ�v����f�x������
���9��X��ۚ���m�#�q���'\9����֠8=:�|��<���7~����4���;��4�?��?o��)f%m�IY:w�(�3j:Vs#VM����F�߹�2�є�������KG��[%O$�w���]k-��P0���
���j&5���� �;ᤖ�xp14�
�bFF�E��TԸ4�O��O���~&�@�@�p���Nk�q(�߶�J���f������E;���bAx4���X�i�H]t���<��Qr�#�K�A�5	��������w���~�����?����K�S*��iY'�����9ٽ����a�했("��rOs���6�Gn�kݽ;P�>�5�����DUtϰ�<@�eA <��jċA��y	q[ x 7j������aG��l��~�fr��4�w�^�R�_���i͍eȽ�������Ȣf�+>����t�jN�vP�Ŕ�İEǄ|�� ��2՟���Q󹧑�4��,�e�8F�4�Ȑ6R���<4f�B���!�.s�����G ����/�Ғc���1>0V����x�:qG�v<�� 	��ul6b� )�����ީCv�"�l�ߘ  ~ʻ�1���^}7�19'AY`�U�@t�\��d�!�|��w,S��\jr3��t���u2��Y�o�3��/�� 1�~���^������ ݶOp��xgtown�M8*�o7�G�zFɹ�l �f;*�C���#����>�eQ����B��17�g%�n�so�'�EHl7��t��$����7�a餱�\��\fB��aB�w<�a3�ԈV�9�<��"��1�E��v7X:!���Z�GbÛ���%ݘ�ٱ.06���s�S�����^FE1f�d�b)�S
��/@C���q�w͒��J�»�1,0\K�� ~1�LfW�y��� 'k����d�3o��t��:�lR��S�0'���,1�K%�a#����?��������z����^wa�&�>�w��J�/��Bw��x�1��]�7ˊT��g���g�����w�%��j^��� ��r/�'
1�=�)�c\�3F��YF%ԭ�u�6m�{���[!�#�5^:2U9��s%�ΏԞ3�že ¶sj`ϛ2�uKԚ`>_~��+�4<FM/#C|��}k��e��mb"�����$ţ�{ؖiu�����?#e��/���:���A4M�gU�}��h����3�5h������0�B!��+�����@�ö3x�;�b��h��ۖb�c���}�� x����m��ѓ.<Dmr�8�;X��$n�JD�X�G͠�l��>��lP^NS�I׃�Q��`p_��t�f��zp��C4K ��d-�bH�P�1�GC�D[�[��-l.\-q��$`bu�
�nw1-�=��Ym��g[��ܩ@k�Q�f��iw���s��<���!�u1x��>����Ӄ��6?�aT��}n�V*����i�_��q�#�E���J�vҪ��g�#Z�z��D�tg�*��E��`	��o����A{BG��K��E*p����g|�gM8�\�
k���f��Nx�N�����r]�cn<A�;L����ދ�[̎�����w}������9 �%-�����< �/%���h��?���+_�ʢ��Rq-@��~��=Scs�_k�7=1j+�K�r���d��~���Ƕ2�Ƌ���
��
`��j��<˵����h�]sZ4�/S��� �{���(��gy�����֦2ʡ�`yέ�'����9c�gE) ԰���ӌ�Ur+�?�Ll���m>Ǚ��l2l*��N�U��E��!dFڀ�mԎ���}3]�������Ԍ2�j�M*�:8j��j��1��.)��������F�x&�{��dg������ާ�|��|�ou��e
1�B�X�,i�j~��p�,��j���� M� �C?�C%<��D
3�S���?��'&+�I.����h5��w��.�5��:Zby��?�Utџ�����= ����pˍo���FK���g�9�3�-����V���)�j�L��0I�0.+��>�����2Y�{�[f*I� �IOhp�s3��J��#�����7��lG�-?����׼�5K��Tz���$�E>���b�
m��m��K��xi�Y���+~r="��{ǳ.(tp�4���`��J�7�s�< �����JQ�?���^^Ƽr�L�/����g�'�Ά�g��w<�@�Ώ���7�����*����'xȐ�*���w��;���4���}t�'W,O�TKr܈$��YIY��~�k�,i�vI9\�p�����V�yQ�0�?�5�^ĤP$8�F�q�d��i*譺f�}�l�xUƁ�pnJXg�7&ΝP�Ƕu�:�y'	tL���	��.�i��iZ�e�#ڌE���T�Q;�ְ�KL��{<�[) ��Ǳҡ*����^F���3��+��F�ʚe��D�v�],/�;�|6o{p$	bV�B�������i�����?�3������0�LWE g'?\ +�8mM�7�́�F��1:�t��y���=�I��a�mh�ĴP��輈�y�c���%h���+�2_�K�`1���G��iz�F^*��c_��p��w=o��%�2g{�U��YD��@ƕcV�ؕ�BVQ(�~�v�"�P;M�0��a��t��r����n�\f;�FX9?�#?��Ji)��:pI2L�V	�i��*��H��b�p�n@��P���Ң�br��Rk5ᲂ�g���U��'�������_�P���P�`i9�\�T^���2��5Ip'�k1>��P{p��1=���P���0��h���6�`�4�u��VJ`t�`;4�v��zƢ��h{��}�"F٠�>zTz3���db��n�i�7�V�!�b�!�����k�.�L�̶\�ӆN���r�]@�	�x31�	Ř�B2�`���w9���y����`&�P@m �$�[�p�EN���#���a�o��9���7\.r\��W�W˸�^
T�b����厵��� l��.#��;�]�c��e��y�}�����>�++�����e/{�T*��@+f�#�5	-�jD4*�5M��#�w������YrţXƲ!���@j�\S����'��m��?��&R�?��m9���<�v(WIŴ�a�ʦ]�UTø���7:R؇�rM��x`GM���M�0T�,��5�=���Ti��J{���&0ƨ+�1� �L@��z�s�*mRJD�L��ա���=���y�UϙV���z��h�EΒ���������^�e,o0j���Z�]�\kP��0���;w}�8��Y~�t��MтKxǨo�v�.+&B!Z.��I%�C��$�����,�+\H4�����E����y�M��AZ���k��f�[��҇�;)tA���i-��I���P����n 1�;]��d�,
1Q�<�9�z�C��@It`M4J���I�i�w�.f;��Ш5a�n�!:�se\i�}e�{��P����Y�6��&xL:�,���P�K>O�}���j�h�W��ssFDʂ�c��]ES\6�՚�����3ӄ��p���3���W��ʈ��s2c�3Q��Q{GjJ���Y��*|��M����琚�����UERyO�,������W�m@�O4_�MF�a�؋�D�Mmap�Z@֬~:I�^s���r׃�����Lh<9 ���@,�cxʺ�آq.�!6���>a���b�y�ա�X��N�^�>Ԫ�k��$�/�|�ŐI7/��6r�Ӿ�p�G[�|T�cvx�2�}�G�N�p��ֆ}������ߝ&m����;A;�]���7�H��5��^�]Ԑ�� 컬Ɩ ��S��[)����T) `�A)(O���ݖ9��Ox��ؾm��Eu��;��5�ub��2���;F��
E��ǭd��4G�z4�A�6v���vz�����]c��!"�-������_������DD�������DN��vI��(���J9���c�t�[-z��i��@� �7�םE�b���,i(5d;_��E�>L��:�Nt}
P�������n�?�9}bF��`::-ƣ��8�BS�`��{��y��OV����5̪y{-�L��_�М��:7�`x��]����&�f�qK6��k9p\�LS���˘�����s�H����0�����8w�ü�>�m�'_,�Ej�#�k��r�X����/[zxe4d۝Oh_i�:6�󜩮NNk	g(�f���]���4|Q-"'�I��z���8�?]�y��U�g���}e���6��� �S>��T�ѡej4
c�N	������ͱ�bg��eb���ye=�G��e��KIj�Y��Q�����V���gu(c.5r�F|9�etD�\��2�@O�i3�ޖ���%O��h��q��C��@Q4͐�Ԇ��o4oz�p^��#��Ϛ���y�� ���i�4��K��K�c5wK��S�`�������\��2�����bD�h��|&�F�  ����ʙv�K�#�A�I5O���%��s;~�0�q
�X3ƒ�ZL����bG��[�8VoV�<��c�;q(�����G�;��lMO{�\Zne�|ѓ<מ��6"W��I�ϲ�O��
7.�b���b��ˣ�~�i��Ѱ��臅9n�,5�a�m�.� \��aw�r���e��K9��n�䖘�8w�-)��I�֤SՍi[+ֹ����\��px��"��H� �n%�'��Lx�O+[ >*�Y��{���;� �Q�[��i����� d?�ղAT�tzѧZ�n��δ[!��!7"M��,؃�1���5�1��\k$�&b>hz�=n]�M6P6��D�"�^�,<}�dE�-o�Š�6�C���D%Tl�GD�FC��v	�}a���ۅm3�I'̇�����/'��B����$B�\��E�d}zɉd�~q�p���=�p�kE^��o��>���br͛>��p���b;�|2� 6����@�����������PD��!�v�����-�(��89�R���;u �R�����ùA��C��b'�\���4�hy'{�2jkz?3�z�j�E�[T�#��Eq�M�}�F�ѣ��0���Y�}�B�y�_Fß��S�-���:= ��5`�~���.�ğ]���xt�˄:ᤗ�#��0~�>����E�r�3���$9ae�o.�KI����n`�������Ҍ���Ck9�"�5zo�Ծ �D�Q	�BU���tgֵqLn��l���b�"�f�+�#��!�����q���06�Ś$r�ir���p���^ic�ϫ�,��y���5�d�<i�����}P
�+�޴_P�r����;ݻ�'���-�佾p�Z��� 0���$�� ��|?n�3 ��T�m�v�9�>�P}gҗ�$�����C�4�A�b�E� &���N��?G����wfJ�����H���=�f�<~����3�K��>w���,��E� ��O���L:�c����\�f�p�s�#<�� ba��n7�`cD����y�~�ﵵ[w9i��]>���Z�����T�<��r|��i!��>��n�	��^�e�|���yNrKZ�A���dY��6\�Or��4f�
�6bC��i/��ݝQ��b��w�"���?���w�u����'�3k^��Oo����ь�ԁ���p�0�@������=�KʳsQ6l�qGjMFG̗��)Q�W������/��Z�?|w��������,?������I��䈗V:F3�z2�u�s§s�<��wy��Z�~!��	��K��i{��/�}�jR�s7'�׺�%�!�Y�s�c	8�6|�½���IVpN���g_�&w�?�2+��"��$%j-T�uP)i8-��VM%N�M
"���m���ȉ <ߝ��	�1�o�C�Iz_Xo��v��m�Iǭ��Q�� ��: �
#y�cް��n4��N�8�s�\{��������']m���4�Ϛ��^�	�V�\����i���v��� O�uϸ�(�1!o	��.�Z�?$34��QҔ��4�����f1n�=6o����������h~Os��f�kÇo,9��l��� �@�X��Vk	�Y$E�:'�13��u�F���@.ԙݥFc���,j�	�j�����#�}e;Y�H:0����ZD�]�<�@&���t��/J�┅Z�BI�vͬ��\H|9Fe�s�1}&u�d�Ny��o���8!`6#'w4�!�)�|n��q������C0o4و	���`^���5���;�+��i�;�=�u <jw�G��7����o����G3��x�B�̺�8�+�;�3��<�#��֯Q�yo�1�='<ҟKi��W���qs}�j���,?�9���^�����Y?!M��:����	~5P����?3lP�H�tq�>Qs��djvu��<��J�El�s'H:�k�C���j�ׅlՂ��B���Ͽl˚]v�Q�~�����ĢTH�����\��K��9?Wj�w�B��4rr)˝���˻��VM�H��M �)���~q��d2e������}�}����
�ģ^����op��Bmt`�N̄�=>lf�Ǔ��mv�����G�R+�x1���f���
��;K�[,�s�{�f�=;��w�i����'�&��u��i�Bi��Y������8ps��䲉�����f� ��[J��Y���L�o|�hC��vI߇��{�+MZ�	5/�B�8 "��\�l�Զ��_��"Y�~��h��
㣎�Jg3�vG��K��M��']QYb��E�1�]�m�сK�7����M�aP���o����(�8�(��!	��,6y�^�]��i�;AH�k#S����D5L�;E��ܝ�N�j~v�Z�쀁Jڤ��N��G�C��I�7��l�[hD���yoëa^�O�JUƄ���3�#�ݻ�v�ּ[�g���M:�e��B�Lk0犝INZE
iS�\���F�Ms�|�n��H�I�$i 5�z�y-a?�HB��%��\���+;�����.�%�8�|������9fy��M�q�9�.�i���RY�]��x_����N�����H*��?Z�Z�\�S��R舝����qK��x�����g>�����MG� ��>��>�������	���Ex�z��M��'�w�]5����گ����4�ɚp�{s;'S��` D�:��o�S���v]с!pg�u�2��R�� x��h�B;�Hs���=�Kl_�lT���;*�w���I�N�E����vJ!z��I� s2���}վV��&�hN��$Qp��U�e���,���_u����[m�;��&X�;��L3������,�z7��zK:�8���g�{g�*��R�|�צ���5��`{�Qv����tW�a��S`?���
ճ�/���M�E{r 2�a}��=�䗣�R��偭t�dc0�͢!�E5/F�d@���|��k�v�-��}ٗ5�����R��S>�S������y�4���I�pߑ�i��'�)`6kv�t����$:���������6����N3ݙ���ʼb�K�q�媜7m{_簟sS�B�m�
�/F%�uP�.��,�:��R�S���2���a����i5��&D��I-+��UϷ�=]Xұ�.���;%A�62�$�$���~�Gf昚r}Q�I��#>na8�����pQ�8����He����X��۫�i����2�aB�)�d�L�y>nK����fo:��N;\4����m^���u ���D@��Q��t�uP�	UbB+6p�m�8��������������rr��. �M�m���B�,��Yq��Wq���i�;m�A7�4�����.���%��D�ᜦ�{�-���=M�h�(�[�7���^���34��B�L���g���M�U��i��U��8`O0������o}�Ȫw�%��:�v��V����,���*Kc���m׋��'}?��Ԁ��s�����)��җ����H��,T�wql��
�DBsF�d�$wJ�e��%DGt��|>k�by���^3� Z(+����̔!�A�3�*������AU��N��1Qu��hK/1�x��P���_~SQo���Tۏ��ਜ�j����̫�O�����Ng�����o~�E{���[��:��;P������������%�4U�<`	8���;8������B�4I*ƶ'u�Be����hĀ1��IB�B	g]xNք��j��3�ǣ^�EM�Q��}������=
Ʈ0�4B��3xd�EB�&�AS)�J�~��_] �M���Ƨ1�\f�1u���[��ǻH=AIRnոv�/���7��^���BD��C��98� p��Z�d�ִ�����hJ?�B*��	㬫�
�ˠ#��a��rŸq�F���o��  �8IDAT<�Tf"ځm���0��[���#�#<�+�u�t�����7���s@@������r�g}�g-CI|�4�.#Tf+[�ʭ*��|�(k�����1��~�`8b(���~"�=h8l`�N��p��ɗ�;:s,������I�LZ���7t2j�%=�{�:x �z�]@j;s��Y��Pb��N6VW>��>8����#/~�~��m8�ʩI������l�NK ��(���r��}�k�e���5�w�,�T�����"�YsM}N��3�;P�4_��k ��U�$�����9��\x�p;u�(���7��~�}�'�:�������Yіm(x^�u�4@�W Z�i^�"����%������s�G�u��	��2ƶ������܇�D��bf�z6 _АZ��V
x�N˄��`����%�ŀ�5˥22�c�j ���,
���K��&��ɧ���-/��ݴ�_�E��G�kK\kF+���Z'"y�	�ѐ��Фx��^V��[���Y�X�X����7��7�r��l��9�7���w|�w���/� �@x���%��_���Zǉ-�&�
�%X�ߌ��c��L�87&6�
�������	��S�_�҈W:�,9�ڝ\)���X����I�z�Ь.�+�aŒ�5��h	V+ N��<��f��ߒ�6���[��V�N1�
�{��{
�����/�b�-�jf�~z�DVN3٪�H�6g,�a��>�]{-��gC^f<N�����S��;���N�"܃���馂�1�j�� �4�2�����_����T���%���|��}]��w��$f�[Cs��L-�bH���L��<uH���V�陕����.q�Dc����J��������YW[�P�Lٖ"UcN�0����:8Y�,���>���1[�m'��A�ӄg��br6k��%���],_\�4r��Y�%�=�43���2���46ǲ*q/�l�]����5��R�[�V/�R��W������r�ŰS��o��o]�����I?��?\xa�1�ŐUƳU�bUVf��U0ӿ�gfg���h|�i���|ҩ���4�~�o6_`��?�c�E����T_�H�p��2كP�Cd5����IK�	w�&�U�LIEn��[H���*c*�"wB�me+`���"�o��-�up�8 ��1�82��v-A,q��\�Y�ĲL'g�s��6��������.�H?��фǋ�f��7tܙF�~bfn��d����0�Y��!���;���<�aú�}jv���G�c�
	�:u�2����h8Hub�m�D)����W =�������:�M���`��q ̼c��=��J��
^bG�p�ω�H���ѩ�d>8(qo�A�b�2�#�������.'1 JL���^J_*�T$�1/ $�wӎ�C�')�/zыJb�;�����A��?��%�.k#wJ�F�$y�e��4���
���uի�l�N7�k���ې2/�~��?�ap�}�H9F�Cy��%b�,�Ԁ�^�{qOl��<�E�҇T���9u� <�L
'Oˍy����J�i���������v��� ��FLа� jf�$8Ǒ����庿�+�R���ჸ�O��O���[��vq�����z#�=k�[�\�$%�8��.h�#j�y�o�v�c,`,���H����g^���{�W��������*��C�y��=x�&�3�����Ek£�ɂ�����;�� �GԼ�%/*�����Z�&i$�<��/G�9߬:���9נ���C?�C�Ꮉ> N�Q�Z:��ِ�ŝ!��N���mk.[꺳��1�u���lǭl�v�������5b�`�%m֬�e����峟���(ו�����k<C���!^��6��]<'\d�� z��~�l"�����R��*`4/'��Cb����2��|�;���w��h�hŖ�C�u���3�3���@�u>5��'��� �I��饈N���[�����ϭl�v
 ����D�*�H��IOHk䄶RR�ϠM��Jk4i	�Ȑ�/�!1��#ΝA�l�g�XM�ݖ*���}6� �����/��n�����aš6DF �2 �/�JĊB���x�;�F��I 2��r��gl��w�hq�9Y�5;~�6�񻹘}������s2�7-,���=ϩ��u0V�#�Fw�c�N�,c{�ql�VF�tv��oDQ��qj��o��ͺ�j�uq���V�������}��ssN��E���ķĮ`=
%�ό��1���=
#�FFP�E�"�5�%����e�V6iܿ޼�mo���tB8xV@چ�Ù�j��􆚜D�(������K��`K� br���D��u2����;�7�r��sq�kC���1�.|Zr��c�tp��ǖW>Y쟌2��>5�&��C#mr�U���fƙ�Mnt���Y�ܸ-ʼg�Iw�B-�*�?�����'�z-[���8 L�b�S#���kv�\������:�g�t�u����l����?��#�[���t�E�<^���v�蒇DtX��J��a�!�u�B�X~�Ŀ�:Y��8x�>G�mp���p�R&T`�3:�B��Ӟ����;�io��a���0���$˰
~��c�mM���m�̳�U�;�ᣵ��sX2���(�˦��+RR� 1�Nm��;� ����	��o\Ì��C8���N[@JCw�`6�u6-q�t��6�z]V���	��4_�� R�_~ZH�0���LM
����?��>�Bl(���S ����Ǧ��h���)a���$˪P�	�����:���83N���[��2�O���'_oi��ՒTD����C@�Vn�ASŇ��"���.�ck�Uy��L���n�P�V�����P*�����r���v�1�Yˡ���>�3�Մg�Cs�lO9��sf�������QhN��fϹ���P�P�"�/���Pǝ+:���,j��+�A2�G�2���Ƴ��L��(GԂ�ГRpR&H��jBjdy"OK��vK u�d��mm�Q����8�9�F�d��}�{�of���;��P����Q��,J��q���2����
��#k�Ǔnb�݇�Eg֌8�8�bjV�F�\�n���P	��Eٱ�������F�3w;�l�����d��YR�uPІ,2~����`�@����ȅ���\͊���̫�3��]��'����r�d;ٞ��Z�i�G��s"��a
 �Fm�
�^W�Ns.y�[�;��U���cbP��!���$~^Y�&�|s0T�o���&�/sV�ɲ�R3e9)�Ԩ����N�8�&#�	W�1�.��!��%s�����9x�^�PVQjA�'��馆�3�6k���\�j��EZɶ�|���C���%WK�'��ɬr���K��y�_���r���s|5�#�A)�2!���5	�i�;U����4��R�]�R����Vd�^����m��~��_��(��v�9��`������t*�J(Hy��k�����t�X�����8����U�:	�j�`�8��LS|&)��RMi����F@\)J�E_�E��=���_�Ņ�$�	���>j����ٟ-��'8�������O~�G�p�ܓh�/��/)�d�
R��>[�q<B��ù8���?�G��	M�Yu7�--s������\o��*�-����F�i�;����9��V>Xƨ�C.��'�*0�O.�����$~w^Y��o��4�\��t.�1��̂�h8��p�2����㽒FpM*'c/�(\\��<v���J�p\^���w�� +٠�����Xw�=I��ⳟ\��c�[�1�a����'~∖Hb�ԡ�������<�9��#��ׯ��M�茉��a;��՟g[{~M�&�+fy��A�\��+�ͳr�浪�k9)S���M����k��e˺{��K>0=��<���Ϡp&h�
��L���J�w�Iih=x�4�r˗�����i��} w��2�vff8���q��X0�S��Z�E��aI��ß�q±V1D��c䀴�kh���1�9|�3�9�IH�c�A�A8�>�$�#���	�F�
��!}*z:Jk�RNP�.O�D��l����7�Vk����.����t���'�"��QF� �9R[�~�����{r.&*�I~�~C��ⰽ1w�(ը�q���f1~<K�;mHf�UZA�*�Nz,��m����IL6��	{-�<B]�P}����w�w����k���; �FIIYƃ�gL*ڷ�]2��O��1α�c��ˤ���w����H^���s��+�z-k��p
I-�ּ�9��Ԁ{���y:EM(� �4��Pe�0ǺK,@�Y�ɑ< }ҳ:�QKKm<�ޘ������[�*9λ%��2%Cǵڙf~�������~D� ���G �L�1��G]&�p.�e��yܗ�\Is�9:c�ύ�ВJ�t�j�Y���3lS۳NF��͘�\(<&�U~�S>��o�����Z�����*� K�S����.��v$�Y��EI�Ey������('�geC��s�F�A��	S��4M����-	&���~�`�4�k��s�A���:�z�5�Z�C2��.p�v+o�5��0����ukǩ�K:˱!�����*�z?�,A�E��������V���Nj��LJ���'>m�u/:E�b�7��k�YtrH��>Y6z�2v@���1�N��N��V�:�x���H���Ni =�H��1	�|D+v��jY���I���#��W�hz� �O�x���x����xԴ��2�;O�Im��ԨS�κ"��L�3z^��˒��6+7_W�������]��T�VaIM���*'^Ƹ��k _��%.x���Ό�'�Ho��7������\�O�o���E&c�0�:���8��PA��M�8���G\�8�D��ƩV0��� �1�P���t�5��L���>w,q�z-��'��I��*�OC`�����9�)x^���B�b�j�� �v�SJ �tw�����HW�{�3��g���4�l:�\rK3۹�z��<�ݥ\�l����E����OG�ٸnM��>H�8���`�[x��ɚ�hi��t�|���ef��	�p���s��UrA��v�Zc�T����F�{���fD%q�$@L;F��3� �"'5�V�-����w���^ku��U+���T�L�������2P�E��L�zQ�컼�3�OGlƆƘN�|���ZWY^���w�s���B. 0sE�2��2��4~��Oȅ�~�����N��'�����4���v��ݹ���{��r�nI[p	"�2/d�<WhӌyA��QIM�I�LS����� Nэ/��//�������'b�d]��$�Ok�KG+���ns��}?�>ۛ6��t��-��9�)��Pg��� ��D�	��������` R�/�K�3XX�X�l3\K]��JC$հ�$�w%��ꐷ\ 385�4��G ^e�
����ч����>�<A���@j DRK��p����XJG~Xm��E:-)�ia��-L���_�y$�`������K<<�s�g|�{�S
�[�tM�B��^Q"�S?�So��N_��'`��F��]�\�cn�mG�Ō����W��> 7[6�������/~IE���ښ� ��S����~����J�4 ���w$L)����%��/���{��	�����e�y�M7��r~�Yo�B�/9Ư=�ؒ�-Z�@8If�ġ-�R�Z����'�������>�nU:��j-hS����[/�d�ߵT�.Gj��P"�Y���5��x�L�I*$��y���~~������!iiy���Tº9ʱ�!衇J��ׯ}�k��ء�q
�K�x����QI�^�E|��F�7(@`���������e
A���x9 ���Z�A��r�8�[z�\}����>�SK�#;k��`�g����|тY�ȼa%�;���=/%��r?�Nxӛ�TJ(�n�V'�|_�_P��k
�9��l�U��xܛ�A}Q:ig��r�פ�>��?=R�����se�E�J$��=�yw_ϡk��ng�^fA8��4VDS�v�n���gc@q-��o��� X�TIJ����N�MP^j�`���v|$�'�@�@=��Z�H�@
C�Pm��pN�ǉ�%&A��oy�[�_��_+������%��X+0�(o� ,�E$�0Wğ���^���<P��^h�(��/��pٸ���&P)�1�+l;��M�Ox�S� n�$�x����Լ4{=�>�`���K�����<���/��/��|ei|�C�(���ȁ�N,�!��9�~k;^�nǤCE�L���8�a�����2#�`zd��r� �9��^k�h����\׺��,@[�<��Lzhk7H90��Eӂ3�,=�5�Z��:�2�;�65b?CR�^E{(*�akc�:��������ƨפ}��Ѐ�!N�3�s��{���s?�s��@��uH�� �@�{�mso����ŌfЄ/>:b>oG�Q;�ﴺa�y��>��E����������ұc\�������.Z-ׁw��0s`���W�������������u�5��ۿ��vr=���`�I��1�-�Ef1_,�Y����>��`���W�H��m�sZ¸]ہ����:h�<��a]�WϺ}ķW���x�+
 1���hY*lO��0��p��HWq�5@��K���\����1T/��T��	|x��_]ޑ9��7�qI�!���! �Ջe���i_��_ۼ��/l~��~�Ȃ��8ݠ `����Y U�2$�y(����;�8R�����^�L�I��:��p��Bf�<�'�q����bGs�Q-�FD�G��]�h(�;����
Au�4�4)���q�#��'I�tZ^���[�����ɖ�v��mM��l�hLLV)��t\�Wڅ�-��q�il�[/9�����4]M7	��0�|q�*][��W���	���F�6���^#�?3��Hϫ�jA�q���ь��]7G9������?+`
}/�jz�g�*v�Y�g��B�s��SN���P�xVh���������£#J�·jF�U���"X��qGd ӎ����P�<y9h	���
�'Z N3~%�/��\n��},��8�J���&��`�rq��g�.u0�q�d�����m�3=�I2�����dMm���{�+�fT���ٛ8'�r1��9�%��@���1� J�/�̾7�\^�qa8b��9�~g�U.� �1�>�4���u�k���ƍ�"�	��������jhj��,U�r��bA �Rp��4��d�{�myN~�b�9y/���vHŅ�΀W��^�aT��Թ���xM����vԍ�7�O���%R�/��/����� �أ!;8r[mX�I�ՄՍ�	��c�p��ꒋ1"������t�����!W��˭M��צ]���`�M��}��L+A 6D-���5���9�����x߭�:���e"��$����XT�
C>��`� � ���k��q�5���Z�
�s�I4�S��sƏ�w��~'���m�F�M�彩m̽P��`�u���=$yӥ}�
��O@5�����5�p�C:�td���� ��f�Z9D�ݳ\�&܎ǋŌ������%yHwS��r���ꏨ�f�$�J&�/�@W��x���vN;�ḁϲI���X��$�L��<Y���Y,��4j\�;��_?��hP���$t~~��T�`5�w�����$Ƿ��/����C��U\k��wU0��r��ߌy�_p�������,�c|y�t�^ř �o�����Q�Q$�)���D'�ǻ�.���,�/?mCA�6b�ءu�����}M���IR�`,%��Y+�Q��X0b��3�ɚ𸃠Yߐ��t��/6��4�SK�������CK`��R�v��0� ?9^���gpX�����zQ�Y�<��\�.,.����`)�.L(�52`~+�#u��N4�c�Ɋ���N��ܼ��� �J�;d�QFZ�^��#�d��?F�V�L�b�G 7�%�@��e�C�N�x�Q8(@��M�1�y3yV ؈��`��}w?��:-���W9@ՄYDT�2cϮ��Ԁs2Oǅm.qjM�ǒ�WV��<���e��ڹw��X� �+�����?���\��\���fŦ�����^aޖ`������,׋��]����}D:M�m�6t��5li'ʖ���6ʶC(/(
�UyWw#G��DH����43J&3��Y.|�Id4����^�4�|R�D�Pj��9��h���-�R���f�$�2��:�8(�����k��۾� ��~�����A��$�+��
O:@]��R��`�-�
�]��7:||<�`O��0�:h`�Q��R�e���f���������+��e_�A���(��� `��P3�s>˼yM�;Y䆙���&j�f��r�:<՘�����r+�+iN�4?1�	äo��˘Գ�Z�*mڟ'��B�T��7p?(�l	��?s���� -�3︟<�ڦ�8�7b��!��I�x��Fn�u��E%CF�K^����n��2��cwIg�JMǩH&Xg�"�[Z(����h���2�#�N؆��E01>����_:\4R��d;��A`�[�<�,�#�*�*�i�I=����Ⱥ�C4��PB�<����|6_:�)�����M�IN���{k	l���Em���(c葤ҩ�<I�J�	�1;�8s���"B>ǌ�F�.U�5��\���u��h�@F:��D����9o{��ʻ���>����P2���]��<3eP�W�+��j�$�����g�3��L:�J�?��c�D>���IZp�fzVYi�?�>�-�
���IEh��j�?�L~�!<0Vd��42���nI@�M�G�Nq�����=�@�=C��`�� �3������6�e�7z+�#�8a<耡cے�I���* ��;rHUf(�	[����w3+O��s&���q�Xs���*�������KA�����N\'�$܋g{��87���L�������,�����b�3D��YT�Ѩw��j�b6g�l'��h<-�0�>*3��?��J�����Y� )�j����rMz=��㚬pi�	@\�e/{Y�Q�F��Ȭ�Հ3f�,�W���������P��uO8���(��*���'��i�M[�3DK&)�4<J8�ag�(>g��%�̶�?����1����jق0���6��|��*@�ʔJV��Y;ƨ�\�|דD����zы^TƸad +��Q7Դ��-Fy�y~�s2輇�6-m��E�� '!�p�>r����k�	�%��N��� �>�����q�16.�A�`ry)_F�$7����А�wr�v*�!�y�k��C�;���0��?�S?�ܜ03��(M��e�y��̠2�Î7
BK��� 1aP�`�Y�t[�\Y�	�L^�P1��΅$-!�M�C[�\��Q�I��r[$5W~瘴l��� 67x徆�ɍf0�OJ�N�� ~9eD�.��8� �o��on|��bU�) 	�5�_���F� ^p<ֳ�������Z���%X��y�p�����͞A6J[��R:����L2L�O��Oj^��7ׯ�h>��?[�4���1�P**�����dU�=�Ƥb�����\)%G�Y��%7�xa;T�G�k3���@����9"�nQ��J��7*e�W�ˊ��N�\�5!�Y�G�8,`�NS��K���[���%#�$�o�"B,�W �����sė.�A�2 :��GY�s��	#�1p�`1GTPL쑣U[�Ӥ�zj��=�q���|S���Y  MFYB����u���
j�0������%>ڭ��ƿ뻾���;���e��1�F��rQ����,���r����Fb����5
^i�̦VM\����LZ�����a���d�����B�JY��O�����q`����6��%f���T&~�`��>v�&�⬐�X.iBls�r�i@;�lp}�\[���5��jIj5���8�@|���[��!���B��5r����A�t^�Y.�~�w�c�t�E"ǔ\*���sF$�J{dd��ajZ�|f�7c׹�U�)I�<+`��=�,
�S�V����=`���������u�ٗ���<�=�G#ϑ{?*�M�j��0�'�xtu�����_X^�	~%�Z ���Fc�Γ��@ ��uY�seup
�TMm��1���s@� �^�Z��Y������iz���j�i�aj���).Vj�75b@�j_��4uP'sMMX�~�1�Y_�- ���7���R���&�dn� ��s,�;[j�9�� H�$����AQ@Q�XY2V�_��Hh	C89��uZMe�IV#�|� �r�(��םj�<�s-B]��rĵr6�0���q����9��a�R���RM/�h~���<�h������bL��#Y�So,�Aʳf���������4�\Y�h��O��2����߮�6��(i�;Y��u�����Tn�%��EMg����E��4߭6|�Z`~F)V�m�X�:��R3<����  cq��q�?"˛r� z.�)�����e>����DI�5����\��ID%'��8�����7,'�����gý��wJ��1*-Fx���蘗�U�ח��y�CX��[k%�yoF3t�	�3q%�B��.��8�Y����W�Q_��o}�[�g�z�;%�Y�p��Sǂ�W��;��;CE\��m�d�K�!�J}7�h����!���?�>�1Ъ���-�!x� ߂��K�iMI�S��T�b_e���r,> �հDnnmeqr^�%�|�'�����ź��^�X3�6钌D�8Dʄ��[�%�㴐O9k�q,�<���:�sg񌭷x�A�0Ϩ�F`@�oJO��j����L�B*�=������7��1x;Tt��̧C
s�!ӱ�(A�����6��3�:�ģQ�D�z1��a���d�Ϡ�SNX��n ��q�vЛ�o8��9�,p#�ʨ���q�p�[	w���Ο�{ Tm13��.J-1N�qo|-�`h-�1�8�9f� (f���%c-w~q����_����n��c�z�'	mF���_���/��k[a��q���A8,�:X�?�EF����+�˱�k�$�������x|I!j8�\yv&}��^�sZ��+�������%����-���m9a���@q�M' �j�)ʧ���}�<8�L���Pc�����Lj5�h�	C?p�Zj�m+�c	��Nt���'����ݿ+��$p��4�jpy�:
�I�ǹ"`"����%�u9�,6��kX�Q�Z�>���~��o��r]�b���vQYWV�(Ƴ���F2�X ����S9�����` �)��iY�FP\��Yݝ�c���ɝfہ�������`r,A@U^�%M$�a!�& vb��� ���}�W�t��ۮ��b'Y@�Z�f5�����t&X��N�೚�C��{9RO��Y0�w�&
?L*�+�i�,��:�>S�SMm/�8X:�̮�Tz ��,c�}7��3��g��vN�$�/Ǡ�RF�9XN闬֦��u,�mq�,��s/J�I�A*ù�iھc.��8�xN��N��y� �Ĺ.��nz��>IRz9��,a�������&�ф�����軓%#4L�*9?8q&�+sZ��[�X3��)�#ﵕ��U���p�Ϛ��@k�&�"�R���C�{�/%?�|5O�RƔuX�_��{�Np�P�E�c�C�;D�X�`O��Ys�1��o�[`F?����*`f�|i��'��nV����\VY'��(�ssQƣҿ�ч�H���uWb�b�fQ��j��R#1[��;�ZD������V.Oj�A����c�!�t@��zr��
��HM1��R4�����ȥ��G����s�i��ؤ�q�=�������1ƽ���:M8ۢ�<\���(�~�����*�Z��(e��C��ƹ�dg��]܆9�(N&$'nz�kn�E*M�Ui+�:�A�OXT-5��H�B�֨\p9�T����:,��@̤���\�	��Ka��
�z�9�D6�Y�T�ۈ	�I� ZgY;Bz�{?���=�(-��Ƽ��P����2��q�^����c�&�n��� ��C~M�;�6�E�9�
�#F�j@��A=8�<�֞��VҏwI���-��c�41iUHZ�u�0 9F�u,���Z�TcG�㽾��ݑ[N@�FEj�n��C�{fVYf�%���]8�gH��\f�'�h�7���n.�g�� ������p �5���w; #�N�Bm�d�4�2?�ZH=�:u+�'�8F�'1�>�`� ������4r�[6��u#�w��Aҁ��?������+_j"�[()?ñ�ְP�Mm^P`��z�e(NIH���+�
�Wq��%�h�+5�Kq̝Vj �H�U���� ��Ť�T3�����ñ`VyJsP�N���H�' KG���/^�n����yV�c� sg�?�O���cܬ�5��rH��2�<���&/�q(S��2ؑ?MFk��*,�`|�r"/f�3��EM��#��}�� �`��"߭�b�tC��sn����\�V.WrqK>���2��H�7����ke�ǆ�R֞6�غ���9��v�����@VU�y�ȵ������PM'��s�C�;<6kN��:���JXu�Eʺ{]�p2O��-屲�1w)�d]U3�6	q��r<mb&��5�g�{��I�d�a2�I�)�U�����L��&��ˑ$
?#q���n�Ԥj�Q�5ـ1a�+=���6���ƕ#��qh��,Uh�E�.˙����sezr��Ҏ�t̩A�I���6$�$	������Eh_\4W|�ս
����6�4�ɸ%A�d������ Ð%wp���.��z@Mذd��9 WZ��U$�]}X/}�KK}
��	��Q�p��ʽ�61UD�\���ǥ*0m>��NI��o���/��|�V�c�=L�ɰC��^S.?7�o&��l�1`�	7�x����W�$������L4��*O|����
�l�U�;�l�[��)�Ǜ�f+گގ�	1?2Hm��'Z����~�k���e�;�ȝ5���*�H֡ �~��8���F�P��1@d�7��:/���;e >��3�[R���D��hՀ�:��G>�4qd�L�����_��R���g����4,/kf : 3�ٍM]��/]h<��f�fX 2��u�S+'���h����P���O*{��5ݐ�+]��s�� �i$�kG�O.� 3���Ea���u�+;�ґ=d�x�[����/�r���^��ׅ�$Ȩ]��ec��z�q�wX��k��֯�t���B�!�@�?���`��SǍ��u�Xx��q9���t�w$����K�dD��R�H�wr�逳�+0�u��3N��05A�k�E���o*9�Z�!o\�qc��J�*m�~G��̴h��X���:�d|��D]bv�aAr/F�CF����h�:2"(�Z����Va��#(4�3�E���g6�IJ�~PЄ��O�ce-'|p���C��bC��i�Xn<�	���E�ç��{�!��f��"/(�MU#4ƕdg�׽���m���7ӎ�B����z�j�j_f��~x�x�+W�݌;���f��3lĸj+��+y�ޔmۣ!Grq��j<��I�k���A.F\ۺ���1���ܚP.Y�$(�=���M�w�x,��ϡ{T�=��I;��G�8�������~��e����sj��t3O~������Sk6�LcK�q�x�(�`��;�V�����U�Z.����)�j)��\��I~����!������&Ub�r_+�Y����(�jÙ�9��9��h�`T�Q'ֳ��;��-�OGts����ޛ ݚ������t��!	�$l@.*�6(� �BDEL0�������[7Cݾ7�R�U^��X
j;&�hd0� *�DTEiA���3|�������o�o�=������~N���;�w�g=���4G���p���zsn8F�W��k��?�K(A��X�Y7t�L�=��O.������d�������Jg�@�T0�w�wO�Uy���������'��Ex�x0��d���K�����;��5��N�����e�s���>��W�bȓ����U��f��z����1��l

Q��I��@�Ș�$NA��~-�35�ǲ�����4�=X��]=#��X5'4��Ve�-��1WT�E�u�Y��H55�� (��/(�A��>P4V�Vf��#���ۻ�����\���F��3�)�ڎ)��Iyű�#_��fO^�A�7���V��؊��1l�]+|{���]5ƶ�b7�J����]߮&�����
�-E��*B�΢H;��f��#`r�z���������A�n��Ğ���G
l����,���:LT�Z�(�ۋ
���},�a��� '�,���9�sk��	 *��6M���gx	d?���}'Ha4�Co|��LD��r��,T�"� "�GU�fi[�E� f������e�Ls���-���w����.|��r,fgϻl��EH^\ೡ8�Af .+; ��gb�a�j��;M��	��K_�Ҳ8P������9���;4@�Ƚ ����<es�v-^z�$̆vk��\3������U�yl��O�y11�r���b��J�<�iO+*�z���7�,��t������j����z�"J�ű����ѽ�6�s,�@#[S{�^i:��À�.��%���/��0�j+2L���l���,lT;N�=��)@E�u��h�`L'�0��Ƈ�Fd���J�4�\L���	M��/���b�ӱ�=,��o�!� *���Y#�%5q%��Gi�RXr����q�(#ҙ����؏��t�2�r�P��"�ǋE�?�ma�f�/��S����l�rL�*�jM�j��J-s�$�4c�b���Y���ۄWV����䳞�����|�����:|�Cz@>,� A���Z�0P_�Aa"S�=+X�V
M�"��U*�c��(Tā��3)���p���8�m�'kH�����Z1�d��DӪt��չ`m��D�h�n#L���X�H��qW%�}����2OL�}���Mۅ�f|ޮ1n�c�b0�>_ބ BK��.+�ȍ?%~��$���c��Sё����4K�\�	�Z���s�8�M^�M��z1�o��V�	��	p�����s\{�E�
�D���at�&M}B���Q��R�L�{j.�A8͟���*��h�����q��Ak뭀�:?U�VWNs+jB�����<���p���8�`x7yP���v�+�+���EG�h�߻�S��.�t`���p�����k��%ӯ��������ӎ�;s�3�4md�����N ��ԩQ,zv�B4Mc���d�h��plB�9ǋ��mn���ow[��s\��"�[�h���X���7���T��N��b�SV�ct�)ɂ��ղ��(@�����\,f9���{k�P�z~֙�3tK\�g���6^�;}'�d�ۜA�~�`l����9��W���1��M{��z���]d��L2���� �)~�l�y�D;	���Eă�UV$�icU�h��u؉X�AԬv"?����HWAC�M������P��`�9��Ύ[*Mz�8��w�h6�S����6���ȏt��#���R�K�㱪��&B��$�c�H��`Z�k|��O?�я)����G�3���w��	�V���y�4���`�$�D_��ѧL
����3�!U\7.�f�H���q�F��lc"�4�-
�����n
8�4NI�.���~��F,��\�}&����U`:O���D:�;�09�w���Y<�ߐ+h�FY]��-����b�����ћ#�M����Fsթ�J�/�ˆ�A8�0d�Y�B�blN<��AxX&:Bt�Ȥ�qH�
����Y��o,�@��6�;��`:�cJa�6VQ��ɐ����n�v���X�j�B�	��� ��Ƞ�2ݽ��6�K^P�.�BȀ���n�i�;K��RMN�h��Z�g�i�7:22I�K��+_���=�cxG�Y_8��y��w�}�k���'�3�k!;@�P�\h>�}Ӂσ�%��q�]�V��'���:��3g�96���7G��PV����0l�P�����I�]疓8�aVI2X�ϱf:����0
B��;�u��7xn�3z\���H!4�j[e���.s��Y�=��7��Z}��L��|��2���e�l�{��a,�w�Z�?*���U�y-2��^���ٽ��,��DE���U���dY�}���s�}mҪ���~�g�h�|���F�#7�]6?�!@��_�C�r��aH��A �!�-��R�4|-ې�ؤ�L�0��(/�ى�2�'�^���5��/W#+si۲��0P������k�f�'I���Y:��/��0�����ogz�3����"���6�Ӆ	�&�&�D���03Q�N(��wm˽u>�6@������~� Nހ@�?�3?S�Ђ��L�:��� d@��K��<^I�\����F�K?DF������4e���]3ID��?����<��uו�c�E>`�@&������a��)� M���KS��nD���1��ʨ�9*�\Ͷ7�J�'�c*U ;6���������]>���-���(��,�j��ʢ#�Wņs�_���j$�E�μk؍�&�"X����*���1��ܓ�g˶�*}�_�2��q;w�t2�L7�dL��ݰ*�h[�\���X5��`a4"���P��K]LˮwP��E���F�(�(�^��-� ���_��.�i��o~sɠ���^f�M��Yo�vQ��v��?�M~��ʶQ�	�-�0�o��n���ډ�����X��)ҭ�R�@Ⱥ��!%; ��9�/� ����-E���5(;���=(�=���U�h��L0��Ô|�Ȕ夽h�_� ��hpb����#4��H��Ʋ�4Ҍ�=��@''<���U ��(���p=
azR�e�C��W���{��	c�	�z���9 ���E-�23
�N����N��R}+�Vy?*e���y,�	��[y�o4��&̱A<��
z�賙v~�'ծ���F{M�W.O{&�p����;G��_򒗔�#I���
��J�o4��{��.�S3��(�8N���R��a9��ن����k%�l<����`�C��횒2���?H�4�X-0���B�������B蘧V�� ��\�UuI8�įx�+J�Z��܃,6��sMl�fM��g�d��R�T���e��<�����i��-�뭴S��s��h0NW�;n�� .T_���<NQZ�M%�	������d����
c�;�!���U��&ev��?���k�gr�D<���7���\���f����na�<�ϻ�գ�������6����A<&� �Ǥ�Y�E�E6�Y8�M�����"G5fA���Y&�M�RF�)�c��(:�ع��}�|o�">�o� ������S�f�c�MԨ�>��h��r��-S0�{���)LxV�k����*�u�ݍ�zt �T��P�l�"4B�����<k��,B8kxʼzD�CN�ݝ׻ݽL�2���T���.�%]qFB�餃���R�jgdڻ�}����{������S%�����{
�#�����׷��嶟7'����v���+��~�n���"�����#$U�4���Ѱ���D���0���|�)�L�wz�H��KAݠ �j��5@q��F3�<�U��V������=�3�B��I&�B4lL���BK��6i �}S��i�0s�e>����~�b�G�^Ď�G,�� 1�Fަ��o�����^]�e��n��]�J�C�)@e����O��v�Q��ʫGgPro+�$�ێ��(�S�;.��i��e-{��8�����O�Y��/�՞k��2�D3��&v����,��A���pVPf�}��ש�h��qg��eV�jw�I!��f�x�W:��\h��wF,��E�y�����6��5�<��ܡ���%h�nLR��c�U#\���>��	��w�q�c�&�c*g��>Xm����J�i�I;��"4���ͫKt�g>�?�9�
ܜ��e`�D0�v>����ʕ��_��W��=n��꫋�x\Rs�tG�F��%]W�㤌M���z@��5�J�c�C�6��s�E�{Ht��̅ӱ��@�z�T��m�ud��, q^���] 8�{��ģ�a������ݑ]8D��v��6-+#ۅ����e/+�e����E%���!J���[M���S��a�G�Z���1�����\��SI�Y��-����	S�b�5��}a�6Cm�G=��%n���G�:�!�>(�/B�L94ˊ�	"���H���/.i�=&>uEA�T�'F�X�D����b��B���b��R���ksE�zҧ��ʦ��k�v^�7mf��QL��;�%师L�]O&�1� [�Y���A|�pD�����^�c�
�y�!� ��Q(���zU�D�Tl$s��0)�.L��Fq��F1�,N$?�W���V�>چ�=���1�R$��}��G�?�%������kvw� te�\�3Ep"����q�dh��"�R�[��L
%�9�)��r�������X�7��=>򑏔�,jU���U�z���/�ʖH�Kq���:k.B�ƐH �U��y��[� ��S�{��Jb-�=f��� $*��|Ϝ�t���"!� cY+�ۨ@��A|F���r<s�v�2]��y�5��(ؤ����,��M�Bc��_����D*f�c���e)Y�� %� SBa�[@����枤]�<�?�pݤc��6Gee�N��-%yb�D��続�?���.� 0B�,��at����A ����P'&�c�Q\����F3MWۙ�<M![hCU]�]�N�z��C0k�f5�bW���/m}�������B)l�SC����S�0�R�[)��ַ���[��"8���7�s$Z���b^q-�^��W4��?���LJ-�Ë\��o�!��;���M<>�������Y�/��/ԙ6�����ۿ�|�h �gĉfv-u"xVk##{�~]�X����h���g���ݐNw�D�`�@�q|ڝ��I+���Bx@�Q���&�s�O�6��qkY]>��/��-x8:,��
F��3�nR�v�D��M���6��Yp�O�QR�J�!C_L�>���ժ��n.�.�D����t%W}��R�Hdz�k��R�?�)�cjB9���5���(��Nt��f�|��8�����qJY��y��h�F"���\�hv@����|���)�!�)"Rw�ܛ>@���2������E�z�օ����	��Dv�!�耢s#T�5`���?C�l�Q��R	E�ⲫRЮ(%�u��Xcu����&HT%��4�cݞ����!H�ņ�I��G��o��b��ZT]���<P�5�3U9=��t|����"��v^��MӁ�c��^���)8�n��v>� S-t�o���`3��cR�}
��Qȝ!8�H�x�32�4��_CHQ�-t�-���)�W�)�ۍJ��`����h�����o�뻾��0i�*h8ܨ��%s��ұ�9}�s#G �`)���	�J<2�_���Q.����uD.��)��;�wW��JO�����>����ǉ��|i0O�J���5�#��]��0��~闦�`Z0^���A]�� ~ғ�����e�����#�fy�Y�e����<���y�9�	y�Ь~��T��\����'��K�~J6��o,��Ŝ�0��O����
#��bYF�ٽ�mo+�F��s 4�!,�� &:	r;M�鼭�$�W����q�")ʠt"" _f�������E����W�(R(sM^,PԞ�gʫ4:N.��$q�M�m;�:4LIU��ϕ���;褁�(��Ƴ	��0M���5�3�-��=�N�qڮ.��㦋�?���q��(h��;�EW"*�~���A�|��v;,�55ZH�� "~V�[{49��
A�����s�"D�%�a�-��=�g��X� j�̡4�%R�G
մ'_u1��1���_�j�T?P�	j�g�.���!Wڬ��a���bǪf�}t_�e������A����Ԁ&6e&�d���:�B4�ݗ��<Um���&�r5)�Paw��8�.K�b�l%�ˍ&2�Ӆ#�\��ϟ}��jW�h\J�w�!j[$ktk����O��X�+�fP��v��-��l��KA C��^��-37,b�KI_L��]�W��2�%��Ō�v�d�vv��������B=A���v�"h� �xf[iFМ��]��,@�%§>gdM�}ҡ��X�tGw�#g��hj0�]5��l��kj�I�Ţ�1��y�����h�B�`8�ť,����K���N쬧��s"c`u��(��03���:�����/�1<NT�����~�4�t5W%�ۧ�}�E�9zs���7��|)�0i����Jngb�_���6���Rt�]�4ϔ��|'�~���(��b/���rG���6�4a�Ӟ�'�iF�(�t �����^�"��xv���6k�'�%Q���ފ��޽9��"�Xf)�NR��;�	���g�-�� ]�,5̀�&��6;S�+�)�y�ܺ��i���,9�ߏ�v���*�j&�E[�_��[�id�k
_��)��T�S0�7?�"\�s4�n����s��m�o�t%"�p"Z�1�t%��e�>Ʌ� ��h�Vi�Җ���b�j�U#�e���J���,�(9���P�}��"T���lQ�z��E��������4�=}�������v�&2�kߏ)[��L6��!��<��|�WVS�f�-Qs��t�mH�q�/�ڶ3^W3�Ϻh�̣4�@�5_��OZ,�WT)n��q�6�>&�?*�i< �_j�[���ߙ5��VЋ��൬qꠤ�@�D4mx/�;Zd��g��8��g��Y���^S�Y?�(��e�Mڹ4٤-�g�g��يI�?���z��皕U���lm����W����LP�p,�{�>����e։��&e[D0�(������E��ϑ߉^�l��\�����Tצ��Od%�QH;o�
��i�NԘť<5/�R0j�����z{�4Zx=3�fQ �u|'�)��I>���=����{Q~���_.^8#{T���vA�H�[��Wzڋ�9e��B�n�p��z�R
�X(���T-j�!c�ex�� ��n�ݐ�\]�1�M2�� ��|�'���>��ƿm�!��iCS�7�s��u?���S8���A�/��E�6u2ʇ�s�ZX���m�hš���W�Q�G5n���J��r��v{啋���>S�]���9n�	B���N2R��%:�{��˩ۚ�L�C�Q^�k������	`��5���;���9g�f���U)s��Hj��>9��h08}�Hx8,����7L����[ؘ�v�^Yo��<;����J�ꖅ�U?\��xu:"�.Ls�/��m��-J�W`��9	jЫ<��|�(�A��\��������&k�f��j��j�,sRM�A��XMl+��^iphǃ�����N����ś����]^@�����~l,P��]�{������X�
9�,�(���@�xU���Җ��+?�b��Zjx)�Ҷ�ɝB@��e&��Ț���r#%��!�Ŧ(�y��ㇿ/���K�M��a)ۂ�^q�Q�#VVze��7��;U���W}�_o�k;��&ج�.i���$ۇL��C.0,F��6��w�@�E��*`S��d*�tl'����v�ʩ��DE
�p�B@�L�oE6�(�>�������!(0 �ͧ��\�Y⹇��t۰�V~����?�R�����0��֊ݝ�V����F�=��U� �[�M�sͥL���!��妗YQ�1��4�ɳ�δv�e�	XD5*�-j�^���IJ��m�Z�M>��q0o���0m�|��q�k�igتQ�>���"?i����]r	\S�%t����n��6���\!|������ŧ�����`�ln��'ڎm;���}�U͉S��yV��<�9�f�<t.e�O�5m�LΧCefW>�w����&�H�"�v���
X3�,b�03���J�n�"�SX/r�uۇ��b���R�+>��`d�Y2Q����.D�`/��������+��x��;K��,��u��w��޻]�A���ܫ���-2�a�p��=�����j+�vn�N4���#�B�����Љ>3�_��9���=c��
�=��%: �(�+�T@��m���C~OM��E�lw�-��kB���q�N�癙�TP�w�#Jfo��������������<��>�*(mY�X0�w��m�7ƍl��6�Q�_��<�1k�[t<<� _8Q�	a����.#(`�,jz�K�j߻�xgb�U��	��YE�Gu&��QϘB*2}
&'N2,��
��#���
T�B�.
]�*��Q��1��S��~�{��ez��B.l/%R�kʊ�ET���b۝h1�Z}p~��Э�쵼�}��f�s�����M�$x~����Ѣ�m&H�]p7N5�'O7ۣ����[��k>��ϵ���| \��=6��x��V���Xi�<��$66P�q�P"N����3�{�
�ź��l��`'�� IW�RX�9���k��e��A�Tf��o���ϥ�'���Ԗ��0s��6��ŏc�1���񿌜?��~��T�a�i�>��n��{p�w~k\�z��fY�9|�ӓݖ�'.�6P��qX���2��}m)pMiL�����z���m�D�aJ��d*���믟�.�`��&U�e�d:J���aS4��ך�]a;&&��|��3,C�&�'��?���/E�a������l�����Ye>� �F�w�£��o�Fi�y�9gx��XG��h�;c4ǳ=�Y�5�}̣���<Ӝ���f������|��vY�G���k����<�-��ۅ���͕ts~�b���{��8�΢a�x��#�wߗ��Z��@�0ο����h��O�Q����UĘ����}�X5����$+d���2������ȗ*f�����t�97�'�!��[��N�;0��^(��s�1��1�L~��~m��5�����/x��_��_�.|o��Tx��	��w(�A.���XC���:����$�7 �Iz�t�R�m���fj��n��mM����*���vyQ���(�/�R��~��`wh�ߩJa:����#�!9��� 08���9�( �+Ì8a�hv೓���A@�L��炥���h#��>����	R�fҊ��x�ϳe�	߻ןU��M��`� Y_�Ew�B�h�h�qeԎI�]�Ϸm�Ex�9��;����~�X�&�/-/��yT�4W�n5""�'�����>����~\�ܱ}�U�K�PD?#���'~�B9�w���uP��)���.�C�]6~jc���F�}���@Q�����f��1i�E�r'�e��|�3�Yd�;����ۿ���w�/�����R_�
6�Q��� y�<�AQ�S��]�R�����q-�sG�]I��+��3�	l������U$��oM
2��ЎRhhc���F�S:�� ��R�w����=�!�(�e�e��e�P�Iv%��%�禭++Q�7���P6h�E��̕i�Y�U��Z��2��6hW��z�3�'×�3ĉ��]sU���'�5�|Xkm[��^iE�U����볛줟v������jy�-kZ����Ҿ�a1b<W[�^8-�w`E�h��t>��4U�4�i6s.��N��hU��ڝN;�N!�b������W'sn�OĶ��&�;��ֺ���3"@���}��1���d$��Hǝ���h~q~z_��fJ�6#Tv��H�3��#O[n[�>̰���ꇚ��E��Uk̼�J� )&2���k�����!|Q�0=`�0�	"�2���_�I��P�.yL�<2�q�m��O鑌b�8�hXz�N����.���ҟ8i'כ>߰��J�ƈ05�o���$��L�a	^[��V���7�9�(o��֬�֊ѡ]^�Ai'�N�R�BL���s����"�ü�ͻw��-z�}7���X?�A��&�Ź�%��g47�tS�� &���1̽Պ]8�؇i��|�L��ҾX����eqWO6����9���
��z�)�^�$�r���s��PG� _lS\��VɬF%Cw1�/��y�<k����x�.�K{�I��Ьg�eJ�O
�����c43�tǉ�@Л��p,C�G�yI�W���N�a˞8��Rk�j��o����kMo@��N9��|�R
�Y<Q/�)h��Z�5�ݳ�"_��˜�ۜ'���e���_��c��� bh��ԴhLp�y�F���%K�*�5A�#�Y=��w@���	�ֶi騿���J8��r����)��N�C�U���i��A�a�����a�bl�f�m������l���`L�搮����Yh �LM�PD����:��eֽ�����i���f֯{df9h��[e��qZ��>�Zi�ޤ��j:����M����iX5ū5u�y쬿��,�t��� ��E/zQ�z	���# eK���ۈ�S����V�7��SKT �N��W����	���m��6ڝ�{mD�x�4U/8�g���C��ԙ75z� ^�4�{U�/�t�0�N�����jd�Up�Z�}���,4=��௙d����H��5tI�x��X}�.ҽ&�����V�)O�����D�p��¼ԗh�3�r~����y��^�ۼEt���K�*H�-5�8�)�&M	_�5_Ӽ��/-�  b^D��	�_����#������n��פ?'�(iZ��Fo�=�Ӗ{��c����	��1.�	Qgޘ.;�Q����ˈ�!�9Z����f����P�e4O��b�Y���N�E(��e�E��^`�۾���wfo�%�gԢ��T�����7,/2��ʫ!ss�����lM�d�]d��Z4��T�zQ��w�~�Z�C�JS�֏��-�B����w��(ur��~���9S��h�ܹP�����g��&�ű<L�+�}���s7����(-3�߆�X�^��f���?�8�D�؀�|��ߘ#>��UE�'g�X������y��"J�j}�A�<�;o�^��R#�"�g&�C��{�S�ؤ05[n����1KfX�p�����^��V����������fH�ۨ���K�,1�O�� ϲ)׿մ/Mf����z�����"��:l�K�/1�8�	�\��FL�<�D��g����6�/J�Ub��Od�>ZieоW��!j[#�sDz�w� �{P���}u���N�'RP�@)<�	OxBY�f�5�H�
Z,Ę��؂Q-�jA�`�+���v�SK����M��,;aݧyݬv������f\%m�B[��vnvz�6��IXk��m��ˠ�v|G؁����Aqᵂ�x��乊�btI��y�z�f�f�2�s�WW�ټs�^��j��"g�aH�W�V�ٝ�цMK�j��Y�7?ב^�-A_��P;X_/��hF��[��k�hgP�K]����n��������N�ґ����<xE?�яN�T���h��l v�uQY�}��t�����p��k���.2o� �>�'>��0YM���MR=i�Y��@0"ǳ �����$b��}�q��CaWs��ZG۹^��ELX&NТ崇�w���������4=ܭ3������I2�,�h֦��JU��n=��K������,B����nF�ԞX/μ��|s)Q-h�����^�ѵ�^;�D˰Ay��C�E����HL�ٝ!�y�i�R ��[��LQ�ݐ�=$V�v��;"H�'Z(�Ȑ��t�{lF8��7��M���}�ו�A��[��ɟ��TF�j�L�x5S�
]�ߝ�Y���`YQmy5ҬA��"��m_���<ٮ<��q��k�d3ȇ�F�j���|utD��f�H��2��!� S:�2�54�/"S�3�;�b�
�4�X��A�ٸ�����r-�d�Qf%���j2EڊP�Ǆ�/h/��xle,Rz�y7>۾6������2,}ɤ�=��Q]����λJ�Й��������R:mP��JɐM"ن�D1F�8���x` o�dʵ-/�E>W�n?���<ِ�����U^Ÿ�Y���"���k����M�y�{
����y��)r2[sY�h�\��0��3��̴�+�%1�+��υެIgh����xf��E�u�����2��H) $m�ޟ��N]ն_HЗ�X����3( �e�����j�S@%��]]�(+�)���+2��+M>H2]�\|�������䋿��(G�xP(�Zv���(p���I]�9 ��5r G+�Y�r7[&�s����X��s]�|��y�4���l{d�=���n}�G��eә�w˜.E��Z�{w��8q� tn�m��z���N��7�����Qn�4��(�jd�����V��O�������wi��t�V�V�B���|+�g55���u(HL1���� \��1V�Ԅh�*yV��!�3Y["͌������z�)/إb	��h��}�@�� ���y�\uQ}�D��!�.�q�K�Ej3i2��)��W�H�5���T@)� �m�D�(�G[M����N��_��_++*�"H� k�9�yN�Mj���R͟g���Y����Ⓕ�tY�&pPUwl{�^�k��.��R�rR��<�h��dz�5�p���_�+�n=�]���¤��2<�2�^,'Ka����8�����]dW6�;eLh\Vxe|͉íe�r�������M�Hr�X�9��7x������-:͚�FiG�R4�9e��B�ڿ��碑%S}>�Mm�9#R��ѥ�ڛ���"�5�P��ڃ %�־2?WP.H�P�P�Unh�Ȩ�Lh�����G���##��X��j�LS�A�DW�0�Z��&U�\� V>�T���&��*`�O��OM;S��E g�@D���m��Y��L&�h�{�*��".�q�r��$�x�h)LHg��c�J�QSH:I�N.�9�]h{��Y��[��!@���9�i���}�k]�jd|pE��q���cĿ3�)��z�_x�QmW;�+�Π�#��X�{���1�P�k֡�"��p�:s̶["��t5{h*��꼁rA�9D�]���	��^����������� P[��L���vhb��n��g�1���[�ȹ�};�~�GG,�'�������1v���f��Pm�H�,�a�h��a����ud�h��1g�2I��b���� ��i���\]s���Y�G���+�ղ�}:gr��{:F]XH(H�
�<�����a_om�0���ń��.D�����N�s4A�͸�Ψ��Y)���NwS.qÍN`�ž��#�7�C$/U��1�Ij�R�Q�m*D)e��X���s�\�e���^���ҧ /��9�����b߅�g�,�Bʸr�����e1b�	J��T#��o�ʚ	�j9������ZDN�;�>M��Gp��ϊs枳�����!'u2\��$(䤭O(��iO{ZA��z���+��+eP�v�����"��,]�=;�P��D�P)�Dz����<GT�0�ڳ��(;M	N��;�6gU,��ue�e��_
���{��p~���Z|�GeM�h�����[�IGc�:�.�}څ}�Ef��˽
���/e�ܔ��r�M;����B�6��p�N�.�s-CN�Ye{�.��{��N�E�<��gKg|���[%��p��/������r�Y���H$#"DЖ��<��!yuTJ��4�j���R�M�x�����4L롧�*Q�<���D߭˩
��4C;\]DPt\����o
9��5�)�'���Q,ЬP��j��^D�z��hK�p4�v-��
�I�v��L�k���Q;B��H���P��
�,l�ئF�t�jt�n�����-���&��m���λ2�<2�t��h��>z&5��?�-�A���d�	�V�����p�Slė2�����^�M>5N�hj��0�\�S8v	QH�r>A�O��(��U(�춋߻ڂ%����8��TL�:|F;��>�k��v>EE�ڴ���9� ��s��B�y��_�d����V%Ul/͸�֢sk��O5�U<U�o{�ۊ�Fx;6=�ڗ��t��b��	�����g���:���~I���T��ez�#QWmk��� �h�n�����=�jh��`l<�d�L�kT�.x�q�[���k������@a-�^�p8�y��F��C�u,뱆R t
�м�R�L�ؕ�=�G�]>��8�H�D��x�͋_���)OyJq�s?�I�"��L:�dSon���<LԿ������s�S[8u@�fd����P"Vn�=�F����Fꕖ�~��)�)[���
_h?��yt���4N�m���w&;p7:�,ҥ,όZ����[�����y Ӽ���E�%�XcзU��ַ�=X���B@S_BP!�U�.k�祶�5 ��4y֣������R�ⶻok>��6w������Ul>�'٬�Ϫ�:�h�����I5�T�ۢ�v9��J��$����E�y�7)��w���σ}�t5J�t�u����O� �2���1�"{��V�yx�m�]4��}i��j�Ӷ�誨IS'*�*1�S(���^�2J�b~.��Y��B\M��y�Zi��4£�e��Y����2�Nc��[�~6��vK�ܼ�&�M��_p�K�q9�aA�<��z]A�~�|
[Mځ1I�����S����e�i�ά`���#��hsí�R�l�����D8����T���p�ݦ�Xt��6v�N �ź���ric,���܅�b�OA�^�+��f�ʌ���[o4�s�pυ�.�t,�5^|-q�r��dw�@�Z���!�4h##������y������<� ϸ���7*��iW��v��}���-��<��YIw��������OpW�e�?,]�4)�>�É����5��񽴷�����l�w����d��y�(��D���0��Q[v���0��cȘk��m���a��/'�?Zj�Xf�Q���X?Lx0KlV��A���Mx4)��Oa8�3�F��E,8�i�o���qͯ��U�ƌU��+
�Ġ�@9bA۠��ݬ���e�_:�2���zj�I��7��w���dS�f����]F��r�ڬ�+�n�E+Ee�V]Z�;�����-ȳ��kHa�M9ߧ��Aa|�tX��7��㘳��ڂ35�cY��ΰ>� �L��GQ�0��u�	K�LQ�暃N��)�ks��ze:m쾬��ԟ\�ܹ#�,cc?!��(6b=ތ	������'��~�p����3��#��a�'�2S���2� ʪ���'�����[D�c�"[^#�-b5��a͸�	#�<��7M8˦��	SE�Wb�.�8 ����/~�#�����N�$�R�	 �;�9䠂q�����A:
JA��m��2�明<K�@"E�נ�eg�Y�59�FK�#.'��z��)#Q"�6�E��2�3ge���A��I�>�@��d�Q��F³4;�`���s�w\����1��e:�h� �}�0�=Z
s�tJ֛H�|�s҃t_P��*!@��=�n�iɐZ��Y��g8��i�.{!��D�ڈ�,6ߥԤY8�����R����Z$�����dĒ����^��xt�s�q9�"a8�zT�.C�VĂ��fM��`�ti�|�++�e�4=d�nskqw��A��Lz����.{$�l�3��(���YK�e�N]�X�=��=H� ��-k��)3T�4�oC�F mpt��� �G���W����]֮XF2��8m�҃t�R]WSD�,�G��eM�4A̪i�`��^��0dQlw� �(�y�Ö���j5~�#�K��N�3�򸖉%x��u7ǝw
O�@O��-�Q1�1�n��*b�Z�Z,��?큦�&:�Tt%vͦ&+�s���O�B�X���7E��	kvXa�ο�[.����g=�\볟�ly���}��ԧ�xn§���չ��Zͼ~��G���_��e�6�~��X�Q'+�j}A����ig��ǔ�F�pj���Ju2�	[1�0�e]����u���S@]A�߅��~���wwW�L�L��N��v��`K��
���3
����������˱0E���暹����~��C�^L�����^َ�Ҝ#c~��/��	QGR�H���]OO'�&]����~i/�X��)�ԏ|�#�lN8ⴟ���6Ox���}�c�w~s�F������2&��{�W���r_V6d�~�~�,z*�]�X�RO��E���GuD@�-vM4�Lهf�AY;���4#~��`,��a����yO���l/�.6|����y�K_zA�^H��w��쀮V�M��Me�,��q�-6�u�u��L1���C<:�I��")�f 	1��l�����&�Գ�W�Y<\�Gx���!L�!��gU~h�������w�5KU��qYr�@(���-8��)w�6�ߝ�3��c���*Z���,��g��1���?��JSR]�oY�.�ܭ7�??/"3��_7��><�a�5��nj����<7�����٘<�n-��b��\lsOC��eȚg���u��a�������i�^���ovmI�0*C��=���뻦��D�	  ��8��H$��=*r?����]�2!�dr��
=�e��d`�8N
�Da�f���@��x+jy}���+�Nn��/����_�����Yί$c�	'��.�ۏ��$"�V0��\Y�hrh�ews�r�pr��Yu�_}��g?{�N���N�c*J�T����+['���~�Y�A`$�U[��� wa�w�Ff�~��8��b�
(�͢e��V��q8�D��s?�Ð��>5:$N����~N��W�m�|ge=?���^J����C�9����sKV���r3�.�F"}�e�p����	z���wP�{�s]l�hkɷ���P�U�Ml���]��1���D�����`��,b���P�P��-����?��He����-������� ew
8(��JN�܄�3��}��Y^�.H���18�D��#%���z��D�j	)DT�sgm�:n�Fѹ�0��6z>�0�dͣY}4K��f�Ft	�d|<^j�ٮ�C~ss^(5�	G����l����D���D�:��oc��un^+�v��[d�耓���2�L�JS���c-]{g��9T�at��ǧ�`2!�q�bR}��xGE6��N[0�0�Cާ����� Ƴ�Șŏ������|���k�A�v�5�R��9�g�g�3������|ڥc��>�f���O���J��K� �3�Ф �G<��g����~y������s�|����s Pu��ϴ�g���s_Y�v�絉ľR�+�E��F�h�j�-��OԶ�h3��^��q|VD�����s��ۜ�v����{,�Q�1���p����&,RϫW\d΅�E^�d���;��LD*L}򓟜��yԤ�K`1�;����z�.!Z��mևN{���	C "PR��!Pm_��W�sElLZ"@wD8�������"-=����W
�T�^� �DB�ig�G��ɾ�Mܗ��?��?�jg�+�Ȫd�k�����;���R�3�#�+���s�M<�O��2%�c��3f�A�"���[�G�Q���f~�nL�ᗾ���f�����h�pck4?ad⛕f�4���V��±ߞ3��KkG�o��x߰��h&;4􇹡�{뎏N�=�sVBp�"Wk�뮛2h���e3�*C��V����t�pkC21�a��z]�r�Z������Y�&K:��	�E�$t�-�w��%��g�4!dZ���6B�2?��?X���C�6M�lV�cr���?��?l���7��G����YD�=�=9��p�'=�I�����s�."Q���o>m��2�|��6R�xj��4��~��ӟ���ܐX53B4q�9:�k^�{���d����VB��dK������*��3�)Z�&�vv�K�0G.t�~^u�aj�ӄݖmͧ;"��+�&4
�f�����q��^�"������+8e�D�V����Hr?<&2��C�MU��J��Q_;횵�Lov���I�9G�� v�/b|��V��ޞ��t��6����
=�^���1��z�0��8`���3M��D"8�ːp�gد�_;�Db����өC�E�w����ɟ,h�6s���H�tJf	J�r�]�j���U;K�gJ>�\�w�jG���(�:�Mb)Fnm3i\iZ�MEq+x�F�oƂ����u��|��R��C����=�Π�*���_U�z���j!�9�"a�y��;0�,A9w��x]�Ʋ{�Tx�|f�i�4�B��n���&��ϴ��c�� �ڎS����и��+
ә7c7�CS-���&���h$�h�UՇ�8���Y6��]��[��NmNgf�ʛ��ߜW��g	��P�	߳�9:�ϋ�!�	�~�}�N��p�}�!P��ឳ�!d��9�<���u2���
M�sʕhmV�LI�W�0��=o� �����<T� h@���f���:B2p��`QbrY�6�Q�i�L�,�I_�r{�e�i)HLڊ53d���g�`���r���§�6y�g�������l�;�<��7������ʃ5�p�#�򾦨�M�}.�5_�}s���t($� �Q��v��W�:���2Hw8����>lrw�r���� �������nj��,A��9�\���Q��ʛ%���.�!�������jXm���ѿ�g��o����x9l��`9���:�>�Ut��G�gݍ��{N��B�{�Y���i.��I;n�B�Tq_]��}�B�b��3u�^�1�Ye�� �\S;�o��1�����Jm�>��}p�f���N`ϟB.c����p�ĩ��#8���ۮX�G��_��E�m��0���Ɵ'N���:El�z��C�[�Wځ���������O�o6��@H�
(��#���^��gQ
�d�4C̚��T#s���F3��,L��U֪?����xS0�M�߬�����57�!f<�QR��]���&���|� �@�X0��(���-.�i�2t�"K���Zf�5������E?��,�̉y�y��xl�.:(�Nw���vk��lU�MlX��c���5�=(��{?�o�3�><�.`��x`,�/���åJW�g0�H�K�Q`��[����x�rY%+�O�i��N�ɬ����s-��~��2J4m4��`GmT@&�M�B�&�	�̊�j�p1�q��fۛ��\��!�+�k��7��}Ώ��E��������?��D�T�Jy���W6����y �v�)�3��1�:��@�_5�4�0�,X����J�����(�r9
�Y�9☣#���(Q��nc����u�f���$���Ex�&��oW-|j�ϴUVz�?��&4�I57S}s�s��~��e"�ݿ�w2�5g{2 >C�2LG�Fĵ��ZLG�舮j�D��h~�F������ʢ`C ���O�8y.���^N4eg��Z�ǋv��s�S�h?�<J�-��<��գ���?���������FG(|�9���Q���-K)�چY��5A�)B��gj��>Ke2�Dg ���K^��/3�Ĩi�)myQ'"lGC�	�"���U����F�������Yk%iq���-�poT�-�r���������=G�f|h���8�d�X`l^��;�SJ��=7=���f��ZAo�ۋ�&��	��-T�^�{Eo����/=�
*l�L�.{�#p� ߯��B2<�'|*�ʈ�&�Z������o.P��Ԝ�����e�b0N�������O���t�!h�P�i���<�'ٿ��d�x�[���t�ME b>��k�����k^���6�Z�֋�NJy�y@FZ�}����T�1��L�X(k�A�_�ѧ�7���T����˄�t@�2�|�䳎tqBԦBvT�cy���٪� �^�R0#����� �ڼ�v`OA1��>���
C:og06?�W�5~�}�v��?���bC����N�-�$�����P:�r¨T�m�p��۾��u�ٜ�F��o,�h�(�XC��y2����V$l�En�äE��2�H��C�d5�ְ*kB���>�<J3�Q�}`yO�^�	���-��@�@���f����@\s� �T匚�|4�v.�y�.�4M[9����7�&��O��V۝ʱ���s�����#�A �!ad�=Z-6�V5;�z�[� ��I������pТޖ����j����V���V�A�c#p�fפq]�`bׅ��i�Ө�=+M
�����h��*��I��@��G�o��h&���� kRNM@������M�]ǂ�W�����i��N2�j�Ь�DTƣZx��07�
c���|hz���}��i���f����]��a�ɲ8g�	G���?��X^�A���w|�\B�R�m�s��yF��3���:W������3�Z���w  ���,��u�ˌIx����#�mv�X���j��;=�\r�
���b�f�����l�����6����VVWoﭮ���6ۡ���������p������m��j��+��S뽕��5���i�;;��#�7 `�A2��	�l2���5&�G�T_p���*�I
��x�_}\�cQQ��X�t�+���ɿsҙ��9 :P��j�E�u�tMYD����O|b�7�aϹN^�Wۍk[�~��㢌 A00��ء�i|;�n���	������_�*~��#�_d��\� 7�P����r�"�f�X��v1R�b6�Y[3W����Dۘ��&5P�
f}]�އ�%��9��bѝ�H�`^�"��k�g��m�k'��ub����S:<q��m��S_X;ٿc��~��Be{pb�3ē����G�Νy����Sw67?�<zg�������U�Q���';E��q`Pj;Q�l)���t]A1KT����S���*t��,�嗿��͓����0|�[�ZTP.�T�W��_J��I&���,2�yf�!ϯ���'��֎Ό�p1L4g�jީ�6ե��%��Ї�Ї
o��u�+� t��c������O�g�9E�:K�G{Ws�}���'���?}"��'��yâN^��m���  G�\��d�A�ӋBY��P�m=6�����@x�I�Y���w������^�������m���W=䃽S��sW��~����}��Woͺ��7�w��ӟ�X���U���Ǐ���g�~v�̝�\��~�a�!�ع��g�_��Q�dK��yلt�#DE�:�p�Y4H{h�MoFmReco.���;<ݿ�˿\�b��>�,�js����p��F�^R��tX^"�e����?۔��*o�ڋ�~�2��~����0}I\�/��/�=E��vJ��K4~�߂��|�0��
Jx7��E�6��p�s���31Ͼ�[��h� b��)��
��=�s'�o��oO�AF�dx�qҡf1afTI�o��!����k[�'O~~p�C>�y�U�>����g7��I7��|F�י����������?_������o�>�՝�����>��1��Xg�G]�&�A�ƫ��1�9�����_}��W��`l����jm.�����8���>�,�(��o3Ѳ�/�2����p���z�긓>���x�R���ߘ�@r� �qcƯ��l���4f��� �g]5�״�BڬYl�M!���E�"�se֣ a����0��PW�Im��� ��"��	��`Yσ8�<Nx�<�茘Ҟ���<-C�O4�VV7�n���֕y��UyO�a���O���es@������z�?񾇝�����'���yp��ן}�7��5ɬ+�dҍ+�MPڴ�İ��F+Ӻ0�[Y��U���:����Jʤ�;���
�Y�9�<8XP�x�ɬ�ʻ�L8�u/�^���$����\}C��&�B���{�)��Vp���l�"{�bV`)���ؤ&/���3��50�]_d�K��e�R�y�o�PTô��8����!g�S�z�э�ŝPCR�+�^XD��1�e����>���2��S�G�	���˦�&G�.K��y���P[��h�����8��s��݃��������}��s����?�����So��/6���hV������+7��*4h���v5�W���_�����f=,��$ʢ�g�����ZA��ŋ1�:��Q��D�:��^&m$��«�C���6���Ѱ[!L�v�N��2R𤗹F���Y!j�'_���8��Ƣk{l�7Qp-��]��y����1HMH�X��6�d��BH�b%������)�B��O��O�1�
J'S�^)�f����q|�jkj3�A��f�5zh?!`�ۍ �������<K�]����C�e6`nQ ��^.�z�<c��9�6:"i4���������t�ݜ�m�������_y���C?��׿��8�������/~�CkW>���F�ίYkzW�{L�Qz;�����~��8Iz��W�cw���ʇ4ḁ��l'[����؛`2P,�N�y�BF#��UY'�s��ܢz"��&�\��
�+��d.��ȝlf��f	���RsrմL��2��3/{>��
%��k�~��R�ÏV���L����/�2 �dLX�+^���~�Ǧ��2痾���ق�O_�QD�=��y�5Ρ��,��c΢��B�9��w�wO��C.�5�����/�����i�maԻ��	���l������s-�:u⏆W�~���'��/nx���1�-?��}�i�����`�����\��5�vm�[/��j�;�bP�K,�����|Q�e�7n1L�BH�Gm�fM��h�+91����w�|�+���+���#g��.θ��L�]"��Х.d�Ѭ����P-������\HDU�%�	K�"��^\􋠂� 8ٺԾP�����7�\�ז�(��HQkk�ׄ�y���β��"a�-����x�k^S�jS�AHsJ�f@栵34��X���Q��Gl.���j�_Yk�������[}�G�u������1�����������7���w�����7�|F�>ͥCc9ܯ&�pƼZm;��xFab:�TH�1kJ��^W	[�{v6ÄX�l�|�:"s� ʁ	ͱ�`�~��KFcEO[�ahV�X~���c���}�s*���lbR�Ǽkxy��	� ��Ř�)a&~�@��)'��3Q">����j��BV�<@˃�A�%��>�N�����%�A�_���xz5D��i7f2i������훠�᱙#�Q��0Zoz�'ϵ�����?������>��+��k����:�I+۫덆'��z�qt�Q�+��F�J֞� �|�b	�1Y��v�%]�|9k������N�L`������L{��f��]:K4��%P갠K�RŮ�(tXD��<s-�<A���sSP��=Hm��P/Y����wY�s��� m2>�!�KPt�9�O�������p���f��F�)Q�O��@^KM�P66���_���1�>�~�0�ߏ��Go-�-�ڇ��F<�/����=�~ss��7���'����GW��9�[��~�~e�k�hX�hkL� յpxY=M䒔�c t�������EH'w�5��
��|
g�.*�Ӗ�m���1�����.aH�h��P����&lȖ5��:�vQ�)L��&<���}Qɩ����6�%@�
�.��������9>��@����m�s�B����z"�Ed��@ �`$�>,�98��>ۇ��h%�$�����տ�Վ��3X?�?6O�x�'������>��kk�>}�7�����`篍��2
+X�{��E{J��1q6YMlĮ=o+�&ֶ�M���%9X
\���SebtCdtr-�I2�L]�EyH��ѱ�%��`wCxX0x.P�QT����R���j�zm�?�Y%���+�.�c�V,ͺ�ـ���O�I�L� R����wO�]��귄���h��)�G�`d��،E�HF�:7Zլ���|��˽<f�7,2����}��U4e����Y�F�n����룍Sw�_����ɵ?k�c���_���'�|���A���͠z�'���kE��}�c�⢎i }� ����sY��\�A�;�
VO��vf�>�/�o�����ȝ!pȩ*v���\��Q�}XA</�������2+�������&������"�1%���a��ʐ.$D�5Gl�'�$�߬{��?&�5�a�8�ۺ
A`E3�&!��I�hl��qaX��25�,�!�b�@x��n;�����`XP01^�G��&t�q�c���� ������\u��'�z�؂��7���a}�����m��k�VUMV��N769�C$���K���-T���:Hǂ81�����b���$�)�c�Q�Ҹ��yWgse�a�ߨ�˖1u��lzk���IO�hٰ�>�$Fp{\?�2�5�@�'Nxۤ����!?NJ�������ctpZ�ŅqY���^��F0�k8�ue�H�X��E��'�s1,cK袻m��rA�]D����������_�k��5�3]Y7��a�f��7h@�]�ɺ�j���?������X�MVȲx"��{��8������Bxp�Lo��.�������k����$e��++��N�E��~oog��a�h0��������V ����1eƆ�X�(D�M[��ݔS-�z7[B�s3�;2�B��Y���jS���߳��]��\ՙ��q h�:�U;v5Na�=�+�<�XQ���gϻT���?�JAg�%��u��l4H��E�3^,���-��@ծJ;�����,���R܉�Y�0� )���h<n��ŋD�P:ʠ�B��VމYw�E���pXPh'Z  �hX���C�7{�:�4"�D� X���w�I����I��^�J�������-�l�ߺu����DgO��w�ε�{��{)]��:��	1��`�"��&Ӹ����)@a>L
xuq,�P��}3�����L�aT�5�!�,���.����H��:׈̐&"�ﮓ:��tI���sml�81��=�=��y�ѥ �]XV>+�8�9r1�8XȌ�YV���׾p6��q�Oe���-�9��|D'���G>򑢲c�!˫�[A�+���H[Ԋ�%����E��FD<^�f���C�-`Ig�<^��M���nIu�<����\�?4��W�7����^�k.�nN�������B�e�$S�����%h۽1v�3X�����3 Z<��Lm}���3S�r��tҩ���`�d���U�d����@�.��䟌Օ�k>�o*��%�f����T2�jDs)�Y�M�x��������3ĩZW`�"�w�g
/� 3�Q�[�����E`cG~ӛ�T�0�������8�>�M�k�4���j.�>�s��\҃y������C�����u�ڡ�f�����Ͳ��C�{2wj'�QDAkG���W�K��Ѯ��;m�Μ���x�7�AU
�*Lt�9b���d�����ΰ (�h���  �3�|��nGt�(��1�Đ�b��,�D�n�.Ѽ��i�E�h�캚�!9FX��\���\��k���)�J�J)�ٯ<��3jf���������N;���#2US��A��A�8;3B��R��{�w��r���cN^�9�ݐ4CE�.X.4���_�Q
�@�w�K{��q_�s�>H��:s�r�>����oIZB'}���]�Z��8o�oj�mtP^����6gϟk�7w��u��n���X�q!WhQ�L�<�o��Ewjǈ��w��3%�8��f��	nXS^6������4mc��ն��K���ڜD����J��մ��E��T�Q�=��nl�p��U��1�Y��EW��w^�WcsQ,�����k�(��.�FZ��h	(Ζ,Ma\/j�0�9#E���]n���U)����0�n%Ys�*0���67�5����Q��.vd�?�wv'�`�[K��Ɖ�ϱQgF(�\�Ex2�B��PX�nD�N�L<Q���N���zO/z�	���qMuZ�bׂ�5�3��U�\�ḿ�lӌq)�$jS�@��*3~T!�y�ť��86
�T�6@`q=�-�s!y����F�i�{-{�qHZ~Ja�(�d\\d2�85A�a�^�v�<94�qmHm�y�}LܨX�;}<s]��vv���/e�;� �V;�KK��8��Op)�n�C��B2İ�ӻ��n_��t�Wl�ﾲ]OW}��h��zŚ��u�9yb\����얦��k���6�O����Y�r�2�,y��X�tR>�Ne�I�3M��5�)@Rșƪ�
bJ��bemUX�>�̉���&����'�Œ1�
)��M6A�]�KCyF���(o�;�S�)L�\8���9j�>1d�J���|�}��rGp�s��!�O�N?F��8�|��WM=���!&��7�����"�;�`�~��߅�-��Rk�2I|hW��N�-K5�щ���ک՝��lJ!��}u�l�b��=o�����iVڱ�z��f�?.a9n7�_h�����y�U�ze���kǵ%B͑���~��D
�Q��r3BU.��W�WK:�ꠅ��頼_M5�f��~��|�Y�����ɘ0�uT<�H8mԗ2�N��3����i����C�{�!f)D�Eϩ~f�L��-o{�ۚ�����X򥱻����L��@�E�<pw�)of?)�r;yy-#0܆`f?��8=���:��ej�fa��h$�
ND�vk�Ȥ�Y�&ΏI�(uo9��N�ܐ1���՝�W�v6�����W}�E��}L�;mek�-nX'U�K_�vƥ�餭���1�	��i����|3l�J�vONd�	��L[����)%ӊ:-��w�I�'[U�+��Y"0e�E�:Lތ���)��>�L�^tE�])�:�uĀ�a3hG�8�$`{��ҟ�fι!���󬝒�D���~5H�l,zj^�gTK���"&�s׵�Y��t��4��?5O���Y�n۴�-+eN^��n�������9������P<���7޸2��?bo�����G�b8��XN�Tk�V+�W��ca<)�Xl`-���L�� �T�e�E6[3������L�a�rɕ�Fl���TSiY|kR�	�ʐ5ⵄ⥎��t�9!y��+��LB��/��4e9~VJ#L��<��$�m�1m����?���~�2�NH���z}ۇ�i�S"���t��Z�,���0��d�q�K��~����9�1�_γ@�7��	�T_�.�M���y�c�C��o϶�̭O��x�Sox�g�n��G��[n{�`�oX��z��p��S �v��={g0*q#'Z����l6'N��
K:[���n���&		&�� ��E,��'g�&�B�(�(��oJ�0Y��qN��6[���ښ��7(٢.��3.)���:4���������^"�4}1$< ��A#���Fiy����B�*�3�7#���1P�1�����W_����d�l�u�!A�fO���:�Ut-�ʵ��_}�u��a(�Qɳ9ޔpg�:V�(hA/�:n�Ȋc�z�L��k��Z���湝ǯ�{�3������o?��t�����k[i�5+��IWK{�������q����x[txr�9��hΞۜ&R����|`�	�gr�s�A|�63�3@���|O��QM�U�Yq���t���`ڃ���q�v����Xe.�
$���}�R%�!ǖ�s\ja�3[����a��?�X�чSM�EC�|='ۚ��4w�	2"Pڥ=^���w��S�UѪ܍E��-}������ c(�ǟ�n�s��/#���ģ^q�"vX�E,�cBA���KKZ�K��^��8�4�L���7��S����{�I��g����n�����ǭ=�Qͭ�]��u�	+Ý+Vʆ�Â�K�{ㆮ��0��j�`�!���:�ew��1��wu��g�&���2�67�p<dc��Y���r�6+����</�-���٢{��D���y�g���R� ү�ў�����1���@�2ce�~A�6\ZO�Y%b�����{ɧ.�6X��s���cjU9?D�"�j�P+�gN���A$��G�8�wT~�\��Txjrr���>�*j��'{�������Qq�x/K8�joxf��;�y����x{ȁ���D7޸r��_����OY�����!��m����R-Z��C���v�J��F���V�����g>5a�a����0�^��WM�����R.7�j9����ľT�&��ZV�ʭnCi�K��3�A�@��0���,�d�/��,��Җ�,��)��Dڼ3\K�flo��B�q *�%���X�y^�6�ϐ*��M���وP�
CFBh�b7g�0��n��E�Ĝ܇ҕ��sσI�~ꧦ��9A�u&�9/2[�=�m����<ƉyTk
a��}'ьs�����rG��h6Z9vb��Ki� ��Qg8h6Z49��z��]�|ss��w>����^ks�
�}⎧������{�z����ںN�I4�8ך���Ѷg�}��hՉ�v�yc!Dm����)�Rq�\}3��>�^�Bȩ��(Ԋ56��`&���ht�Π���&`V��v>m��q- D��/�lE��_L�h��?j;fF)ty�DN^���A���O��6�'��6��ΩN���H�
��d�M�cY(E�)K����v$1�!\��S ɬQ�T�KH�����nsDQ{�0�uY�uu)`�&�v1�0&V6tN��c�X�O�*��Ѱ���ޠ���������i;u�
�a����gn���S�������7��?>���Z|ݟ~�/����/����x����+(K�&��+po�LG���]��v��y�7壘�D6�3�©�����Pb5k��P*�#/��mͲ���|�̧J)��ȳRHUJ�q��j;�1�-C�,C�	��6�@��E����h��{�Yז��ꈊzLs��̞T���3�*I�1Ρ���uf��c��9W�N����]�]���z׻�Ü���ٮ\�R����	�r�1��t�M�(�u��i�����4j������[]+[����Q;N����͗��h�;9>l��۞������������w����O5G@W��3'N����in��[7��E�v�>����:��~ �����}�mF�gt�T��.�<�Χ?��� TO:�dl(F]T�ļ٤k���0��&`��L~��ɉ�3&��E$'oz��=���p.��E�BB�f9&GL,�:*C�xT&��M��qн��on^��וJr�%���X2Ь?�׹�V���o"<#�����|Ԙ��Z�?�ݖ{���aoeg�26�kK�o�� ���ŃV�g�;E4���#���z�+v��!?�Ʒ�x���=D��k~�M������o���7����ۛW���ۓ@�X�܈�"vx������͸��|�T��F�ZO��R@�z�]�ݵ���|f	���11E�:���oR��!Q�IJ��	�|�/��5�����늶1�Y�1��yη�LEN�./Q�6����}���0��~N�0��-oi��ۿ�b��pNa��w��1�sc>!��(J�v:��6y���< ���
��;->?�vJ��x�L2ϲ1�p����J�P�w{p��w>{s{�����#����_{������������s��So�q�\󹫯��/Y��5w���[�~j�mQ{|����~��/���wƏiGU����Q��\1]���{�ʉb�if�V�J-"m�NLQ����N�����$���[Ln�M|���,^��j֤�oC�f	�㶩gy��\h�q��(�4 �%�[�N܃����#?�=���ȏ�HI�f_<l�V�s�K�dF�8�� �9����.��L��j���7鷝�س���6	�\�l�����R�E��e���(��IY�5��Xȭ�H���P���Z�w�k�޻}EsŽ�w�=����W���˝��w��_���w����o�f�8�~�n����qjcutzx���z���YW�u�3N�{���g�y�����~����vo��=��`���a��P� .	��������6ᬠ� -S�t�
+
ΐ��E�t��愫�&\n|(�y�Wz��&�	�S)��s쑊�&C!�4작���A@3��]��k�p.b���&RDș�,E;y�k����YD_�a��������[+��	�Bg�a:��o��X�|����Ú��,�T�ﶝ�{W#�Q����gvg=럍mV��b#C�#%Ĺ���-nV�H(\r@"6HH�K�,$�	�A � !���(��8��z�;?�U�{U�zjz{v����'��������W��{Մ�q��ѣ���EO��VU�*ݒ\<�[Q@X\۵+���0CceB�W�3$I��Fl�ɭ���R��^>*gO$���hddf�HrE�M.~�o��^�i[�Z�<���e�I����C�4;�,5�'���Q���PF���=�1.h�%�F������zh����XK"&t�@"/���m�_А��2�]Q}�MQGD�D���K/��E�W�ԡI���|$ȓ���(�>}:'�li	+l����Z#	�ॲ������Y,��PG�:]J��K�U�����}��j�zA�H��G����9�`�$�'P">t�P�lI��,(ݢ�IS�lH��Z�u%�S�oBu������ f=[ȹ�S�/|���$���ρ4�'��0f`�`R�TSHÅL�D�Jq����+6� A��D5����cB`�I�U+sY��(�y
ucB��\g�h$u� �WR��P?*�a�@�u��4;��9�� C$	3C��^;���`�Z%��P��,������/�B�Ӊ�}�a�t�~�!_��gb�'$�F3>DqUg��_��A�����&w|����'o"�$9�h�$LsT_Ɂ%D$�^z]�*��"��(Ġ��_v�����Q�#�:}#$e,[tLB{}�b��%�*IȾ�M������E�/LH��.\ )�����bJ2�?n&ѿ�8y<N�Z�
FNC[5-������a(u��E���8��x�ep�U_D�i(�Lڭh7Ƞ�3&l��ք�d�����R�cf�"�����+�2�5;���J���\]F�垅��sd��}�Z�_�����>Ń%�$�~�,|H���r#h#m�&�N��0�=�a��!,w;$5�ݭ6�+vOKܓZ�:$�:zx=P�g%�Ǘ�}&�!����Ɨ:'�Dj؝4���Ȉ$A$Q�u�e��qHڤ�݈o�l���y�}Q�j���^)�|1P�on���߈�I�e�쓳��`t����Ե���$,���|���b���Z��w[O@��Z�yh�PYG�*k5qKP՜%7�&�/�<=l$L f�����%�Ђ���V��q�q�Pd��R�}x��5/H�x��$2�8k��*'����q�U�4v��đ�L7�V$0r��-$�����m�{�( �M5�����L
 M��TK����#�@�
LIe&h�բ(1^�ܶ����F`5;ٮw���}�Ң]�o��ە�k�B���ۤmc�7�� A��oޯG�_~~�?��'�~�����I��\��]�>Eg�S����Aq�A6��<B�R�����?�䓿y��W�R�UIU���O>��w~�R9�Jh4��.JH�>[�\A2t��Z����1�u�"�J�
͜K4��ƨ{�&p��S��њ{i�Φ�i�X��y��u�S6��T��>�|n���k��Xa������_-5��
�@�;���{(�=��r�F+�(6�.L��t|��͕�F�ïK(�I̋1���l��� ᓄOt�ٞn&zIz��z�[��F���|�z��I�4"�dgMs���o=����:���b<~c���v�>�0/���]��X�F��z��'2�2�vY�ב�2�% �,y��ƥ��:�.��y��2��WweŘ����M�Zv~�4e�KR�pz�!cf�f#0���s$L�������Ҷ���TM�r��)aI9S���U��(�߉9�7�@��E+�L���O�E��v��(kk������ҍ^D�Ϟ��Mb��r��e:ύ�|W�2K�A���H��<�*�&���bؿ
D�H��x�g���$���^�9�ƛ���H;m�MYzTe|�F(����d̝����a�bFf���ˉ¦҉��L��W"����N�)Cʖ�P�v)뤬���|�����+��|��׼������n�%�N���&Ν�;/B��N�|?љ�T��0c�����D����̩+� ����H��fLnI��&�Z�� (кo2� a����:�A������,�{���ܢ�����?>��S����떂}�������?|��Q�[z>N���1�b{�*5�!s2��*"R)j�'��b�~��v�Lc]���c���-�9q��'evQ;�w�~��V�LsI��/�'�hێ:��V �$cn:͊v_IG�<���V��� ww��(k$�A����3�aK������0Q�D7C=�τw���|��=�Û	mgV�/H)�LLL�=r��/���9v��ۈ�Bv�ң��S"b��hvi~�j�>[��x��1Wh"2C^��mA��r�1j�ʎs;�k�QG�H�K���F#�褶p�ɮ8�J^H֙�S�Ga��J������LKnE�|�2f�%�F$(�k;�e�ۦ��u��J��󗤺��-��k��i�Ӽ��n,ȵ�����p��E(�k�����b���;�Y�!`#��>�j v��|8ۯ��Q&�o$��h�Qy�x+"7ȹ���Q�V�-�7���ܾ}��<v��^x�O6���[�OO+��'��F-�}�+s_�K��h7�<"d<�2U�*�@sM7\(�y%�:�� �I��u��I�ܑq���KA�+!gn�������a�0k܆�]L�2W�Z/��Z9�K[F�Y� ʮGm��	[� 8|]e��i:�U}�ݟ��M���r���3�C|��Q�r�5�g:�	�`^DѲ��(��qeTF��
ɭ����$���x��M�<@�ve���o�t	ig�.�Yv����B�le/珅�k{֑Վ�g^q�U,4���E�:W\_��5�z��}tٟ�A��Y�.��o��Q���j�\~�#���FGG[��M��?}�����O�����_߿�={���=�3]x�[7��g�V}��lt����X��iV������{Դԉ�d�ⱝòt����p�t�)T1PqUe��E.�a�P�]>�9]h��k�/����IRvS�	\�)��C	Fl4��}���FSm��n�.5,����r v��͐�� �1-@�7����/
	�Ur%��@q���r!��mvg�င���+���(p\d�G"�*V<�Q4�rҍ8m����92r�Y9��t<����y�N�8�nvS;�l]�#|����,;?x�F�V�یu�a�y���=����x	ҫ�j��c�=V�8r !G%�T$�2���E\D:DR�}^�х��l��,�����7H�������;S>*��r�A�%��|W�D����D��D�8�@����^x�"�v�DĘW�	Mb@�}�����d���Í�{n�̙3l��>�R���f�:���7>UK㥆N�D'�v3*V:IAք&E��ɉ�<�D�I�0�x9j�Q��	���$uǪ�y�J����ߝ9>=���٩)�N�T��s��_a��W���T~�����ۋ���v��N��u��g�u���Y�_��SǻuuvV�LN�=V�KH��5���|���LMIv�<:=][����L��Z;Sz)br9fzeX�>���
i�d/٘�Sc�gV�G��2�>g�k$�s�ߥ\Xے�8M!���Gؿh;� a?�}��ӄNT���+�J�b8�D������_����x��x��ָ�����C�ML�����Ǒ,�-c��Eh7@�}�СCOMM̓���AE��y7HV��z��M
RfN��Q�^�a���9�_fl�������M�k6��l�������~���͙����by�w�N�=i٨2]��S�ɖ��,�-���I��2�!&3���]#��X�ZjT�� ���Qm��e5��"������A�w�n���V�&z?������20��(����k�g��Z���R%�@����Oq�ʝ8��@r���
�U����0^,I_(��r6 �
��Iv�����;w�Lϟ?��8q������4<��U���v�h6Z���.^�����{wף�0ȵ�H�E%��@0�SβD#Y%ZF�8 	��L'@2F���r�w�Q���Z����DfQǑ�*"IϦ�OQT�<C:��O
�Y����R)k'i�J�T"ɡd�h4�������������{�l	oA=s����W���.�-����إ��y%޶��l~����6ν��<y�d>�1	�t�Az�F �-�	V?�kl�0ξue���NS���N׽�� �7`+ ���V��V�]�q������e�!k ����v��Į�I�ㅙ[���/�����!��������GD��F���w���p0�UL��:�;I���ή
׶/r�'��ga�dgaa�llafbbj�p8�R��hN��҄��


	*2.,B|J�?���m�X0g�?x����sJh PK   c�X��{	  -  /   images/62a7f633-b11c-4122-8d1f-7a295c29ca39.png�XwXSM�MD��DJ("���"�H!b�RBo
W� ���D�	(H��"DA�J/�K(	����~������?;�s��3�wΜ��sga|F��w/�����1a���t=K��a�R��6=����,����D4 0�k�Ƈ�y[��aaޞ^�Uꒂ���TwH����m�����$�?�3M����s�C�G��j��j6.���رc��+iJBg�޾/���%f�jO���R�^1�:�$A���)���V�n!�C�ip�2L{[T������ktdP���j.���}��z��������U���x&�R���7���ae�>E[,~_��q7�L�5M�((�l�x��T/~��r���Ou�	b-�䶅T}������'�[�8TW�X�����k`r�ȵrq����=%�s��W>w�_����stt�r1:��3���VJM��0+ӎ���������=ƞ(��=��[�p��[%�W<P�3��sQ^ieG[�y�VX���V�ݩ��H�g\�맕��R����|�t����9���0���X��x�Y�`0|Bk�����bj�kixG �+��/9(�{b��Q(�ӎ���+v����CCb��,!�b�!a�j�h������p.��)!ؕ�n/i�ı�;�ډ��y��5$���c�k�X	�? ����^�Y�i�����	���bj�
�_rPW�SVTV�*)c�T啕pʪ8%U�?�k<o{G����?Gciξ��8,6  @!@E���URWW�**c���Yy� _�@y��t|�.��.D�5����WCB��$�=�r����B��h�URP�����y�y��1�=����������*���t&�}�����^�� �H�y,���}|O���s��i��������Mp8��
Sr�����`�K�6%�~���wLb�*
�b��.k=2���A��hH��,��"��b�t���S>,�x���7�!���1�?CY�U�))��E{;_��lO�9���XSvq�sr�zz8I����8m�ћ5�?\��=||�<�:�{�"�^��N�E8E;%���T���Ԕ���j�Cj��TT~��	~k��mo��7�va�.;���ڞ�Ó��+]A2���ן����<�����!A�#K�v���+�7� g����|���v�ǝX��_
�
��3���$���ow�����u���U�<X�˛U����`���q��Ω�����\�mt������F}���/~,\X~3��hr�פ)g��:<�!9��q�����+��<g]#z�P�'I�Mt�O ��r�U�,���N��[0�^sz�L'c��9�ws3g������ژ�6�(}#��a�.�����m��Q�g� �2/�A��+��z��[H�=�"#NGH,�����c�_��֑�L�;��/j>����^,i�dߛ3�Z��$O�9WWq�� �/�����ad�S���A/7�
64��E��?�=��E�y�3���)!�>Su2�u�����@�f����4�k����H�{θI?�A�̟aQ��	�6X6�ڸ���"W�]�?T��f<5.�}'~���k�Z	��P��ظj/ЄRo�E't~�FS`�|��O����K�h��S6d�ʢ��&����e�t���&���˗��Zd��~�a�͝��K�P#�ENC�V��Cd���;��� ]�7�vrx����Y�{����~:� }LN1���KZvrP�Jo�Փe��]����ʏ�ކ4���5�З�N7�[���2F����B;Q��@=Ѓ?�>�b�"��l�L@�h�M��\�-c��^a��嚂s;���y����3�,V}���j�.�df�>���[���F!md�+�^��q�������,�/�h3�d�x����߻-�^Eӣr�3i#�Q���A]#�<~�#sq%qr�S9]�=�˅��m��e)	^�+�~eDL���U�Nh3��p=0�h���<�<��pD`��+�-'��Fg�0���G�,t��� �V����1���V$�<�����t���b��5Jf_�\ӣ��zRZAn���
�e����&��x�����O��Y�9�F��wߑ?Q�>5�5�׌3��>6o�eL"nm-:g��2ѣ���O��$������gg%%��U�^P���8B-�,mH#Z�8��$�
b�}�go�g{��Et�/�A^c��������kg��Er;��U��	���j୽ɓ�iVV�]$��C̷oA�C���l=Z�8.
>�N�Ș8���9�ԏ��l�QF?5[*5t�j�B������mȝW�����F��?	<���g�|�Y95$����9��%�A2L���IM��J����;�E� ]�+I�M��F��l��2��+�1g8�a��+�g���Lzx�g���4o��|z�)bq�ˎ� ��>��n�\E�[m��"d�4zr�k��W�������
^��X�!՛���EUbԕP�̳�����k1Uy���W:���*σG�c���W���gF�_��8j2��`�����o�{A��"tӗ������uÝg��p��$�=���JN��7�`y��JLoƍ�s�S{�w��������V��;��C	c���N(I�+m�	�9���;�7�%�]M�OM��;t�y��*�u����1@�iS�yT��f.�@h����fY��$%߈�&ײ��Z���������6a�W�� 9��l�1]"]c��,�?j�#r]ԪiuOV��Q؜a�*������U�7=�C�;�b���e�I�'Б�tkZ޷3���Ei��H�ڞ�u$;�h&��ǉE�gUT*���Ǉ_l�iVh��AnE�#A�3P�NZ��l���	����oF-N���yC�v?�5ߴS�Eƒ	��ӷ�ْ�ZV.�[�Q����V�}�ܛ�{&vv�A�C����o�A�BY�Z���s> �R>�2c3g��<�"��V�׭�y���e�`�AM�5�x=:�L�L�4�4�>�=E�u_ Z,��Z]l$����0w�(-���1��-X�mkWQ��T�s���eXDm{��^(ѾVQ��R��	c��S`b�*N%J��ݿ9YO�й�όb�eO�\���ba���Vd �k�%s�{3c?��^n�]+� �l����Yn�����n���Fjh�ٷҏS�����0�O��T9�@M}K���%㴞h��,G��F	wT�x��Ǉ2~!F:�F�s�ř%����`�'�W�~+;_�d2!��e��h�eV���@�@ޡՋ� l&�޳5�@��IHg����o���^�2L�9��*��8�6T�(;������ 1��a�5Ő;�y �	��h4πg?x����[?ؗKSIK�gP�+ǅ�^"{�uE��p.oN���p�5������04�32��?�/bP�ka�W�0�?�~r3���\%j��m8�ِ���Z�8����Ѽ�}[�Ե@Z����`�ٰ,��d�xDï^�W-Y����=��o��bn�բ	Qݠ�ˇ�R;ܭ�:(�L�3j����O��\ [��*Ћfx"���(LPa�#�"兏��-�Z`��կ��(��"��4�q�'l3�bJ/��V *:�sS��hō����|e�S
:�gO'��HG�;�h`U��J��Z:3A�2A�ܘ��{+�]�#�e�BْFԙAhf7z���ɽWS���N2�:��}�&�!����������7A������>�hMT�#�q3F�[;��#��6�ѠR�}�i�d3�r7ڙ�C����G���y�ҋ�$Ԣ����h�_���{wυ>N[4��h�Y�#�.p{��D[��<��eBg{�" � =�`n�k	�4b3
��P����}��	/$�|���PJ��]���F�����
(5|�<�i6��;}�=3$��ϵ�Ȇ���vd��S�����!��O��ڱ�k��޽ �-%_�G]r�l����\ۇ�l��'vj�b\�1c��gD�o+��B����F�i��F#�(���;�%CiD!�)2��t�[s[�:��ī��NoKY���2o�#�B9��6
�W%c�������\d�t9Y�c�(J���UZCsz$P�|F�{���ާ>�¬�(p�CGO[���>(=�NO�7-��_�i���6H�z��\�N�Ci-���io�ѠOp��Ew*�c�;d�	�q�����
~_��SΖzx��z�z�K{����� X�e0��<��U�,ު�����f�����n>�GL�T�5��6�=��E.k�OC��6G�(Ti|�朲$:��t+X�����.|d�����;�W!��`>bys[#^�te�V+W�Ɔ�ud�o+�(G)��~IN�!TF �[�G�R�/�W����Z���%�Z�7��(�m�v���9���co�3A�s��qp����D��6�[�@��P��=J{r^��[�V��u��	j%r�P���u����|w7�J8ol�f�N�R�<�-���`�Vж����_N�	�Ol?z��JX���!`�N����� 5e���xb�����@τ���
��Y��i�'9a)��@�� ���HU-%���=��v?��=�6�@��U�\������Z�˿r?�b㧚����_yua-��S���l�Cg7RZ����U�Bؔ�EV�e���ݛ�>co���ߔ��y�.��\�8m,�灣[���UY���UµWJC+):��6�^�s�,��D��xy��꼰0�j�U\�[�J3�jTy'��}��p�yk�0	��Z�ƺ_�h������D"�H��r��@�-����O6ǥC�j
�Q`Uv712S>��6��u����rӄ������[��N�����ɈBԕ���Z¨����v�7d�_V��.`t���+��p]d�A��D�lEy����T���f�����a�G�w{z���J�r}wF�(Y�æ6Cl�S�m����G�����:��ʬ�n�Z��2i�Y56Y�/,�6~sv2�>+ݻB���ƭ�+V�U5�Xy�!���t���<�m���f�ۋ77X����@D�u�۔�G����<zE%q/㗇}�n�L�:{���i�).�)o-	����Hڅ�����QP�:p����(������ ����^߅��zC��1��@����,ΑBA�����t&��C&Q�_���	�-�`*�����/����]�����l�����W8�2X������^fձ�o/��ϷA�2p�ܣ��$�c��~�E�k.,����_�z%ո^D�W�o�	����`��)}�6~�g�d|ʖ�tHd�L?�������d����se��f����=���XZulf�y���׷<��sy����y��;�9Î�ս���~��}�;���=�U��Z��9�U��3u�c�`э-0�W�)�gCL�����=euP���<� ⎸E��U�q+��i�s���LʠM�l~`{ٰ��kQ`,�=�j�I��X8�����#��]�Zt?P�Nk������b��
Z��Oh-� W ���s5��kb��wC���|c��򹎼Z���������n��~�D���;��W���޶Mˋ�����P%;s�^�y�u��(�2Y�U�����dY\Y�ǧ�ǥ���<�z�ބ�Y�<BˢcWP��#ܛ{k-?RA9�u����	_��3ђb��E����E4���.����Lj�'x�$� ��E��3O���}y�����'���j]�7PK   �b�Xk���  ��  /   images/7b670e17-d5f7-4cb4-b95e-fc2ea835e4f5.png<�s`���>������mc]�ն��mc5׭���Nm[���x����}�H��s�s����U�2  @���P `!�3Dx�'���Z�_H�2:� @b��T*��C"7Im75'K7��7 d�q�s53q�`q�f�}.� ���S��9]z�̷�^^d�ϔ��1�W���쳐��d���)�������<�������X_�~�~u���Z�A�`���<g��6D�cl���?�@d�ݕ/�`\����Q���D��?$��7H?����ԇ��VF��x=���.���=s��K�������C�B /�v ��'����vd`���Zf�#�]�+��%�D9���p��[!�|Ə�AX�Ti}��2�UvG���R�C��)��D�.��P��M#}E�w��TG��l��#����af��b�fo��FR$c�qd$qd�h��Y��!�a��)�/�7*�v�n�0w*�fx>#G?f��� O_����A�Ÿ,cw�3g�#q<��g?컹"'�,!́E���y C8#Y?�~�1#Q;2$�e�2S���H.�$�y�T�＃�2!���j�����ݓ�p���������C�%��b��gL��"m�A�٧t����!��<x��J��w:J%������8)[%J�^fJT������^n¼Ā3���U{���r菮�`�,��w�͖�}���B����_�1�f=���ZORg��Ï���Z_��g	{K�򹗮�%y6ʇ���m���d������+p����=�7�U*Zf����.����vN�I��QN��(;i���S�~���2�c�9��8���MB�g�)�X��8��H__��L�9*PyB�F%��cH��F�m4s��ta�lr-e9�&�_"���u�+�4�zy!�<�E�W�@���)s��}�6�J��*�ߟ��!�߁�\�������Mc:���W�3�%���:��H47Ҁ�r�����"��<Y��u��N�;�t���|���lj��!��R��7�dq���\5W��%��$ R�8�������P�4;g��V�ߌ�"����;�����e=�r�����6�G&/���7a���^�ky�3D{�%E~�"m=Č�� ���;9��+M�1�o$�q���m:�l�_/�Bq��������f��w��Č2��ƞ������.�,���yaR͊��k�`���%��{� d��ۯ@nҤ�ݍ#�b���#M�C~EO�}�\)ȣ� s����qJ���h٤�}p��#��X�O�Bѕ��ô�o��5l<�'�OU���o�o,\�����xXn������oɓ]i�جPX�t��Z��m��>�����mo��EJ�tV������)d`H>V�?��e�������J�F�R�`�Wv�|!�eu� �/�E�����?��'6#��f�=G�A� <�B��{rQǆ�u�S��BP#�H�L=�oz ��W�y"[��/&��/˞��_��nB盥���a�_�P+"l�HJ�||��ԥ��Y��l�s��씝��̐U���>ets(����-��g�s
�����7��fi�Φ>���G������G���7�c����*�jVj/�D�.9W6�h�؁]i?�/�+@h_��8��ؾ�0˅U����ݐ��s(�bZ�e	ښaF�i�S;�,���U���E�J�Z�+�f�Q��fX�A'���83t��:Gg�!�;(�݈��-����G�O7��{�pؓ�q��sp��o�[t��q�-g\5�#@���E��nqg��g��Ϯ�eM'�o���՞(P�ol���r��f�Z�e�Z�W�#/G/v�N>ą�A�<������I&',�-�>�l���<ɋ7�6���4��'{<�Jc'��И�����D�i���y�-���������ǟ O���o���_�7�D>ܟg �Z��H�y�|�7W��+e lw36�J.ح�*T���Y5�?׷,��`��к���O�� ��Ric:^��|�;1�}`�ޓ@�jb#@��<��G"�(��'k�ᖫ9��/ ?xf�41ũ�J��툌D��en�1�2��AvFoG��LnҮ��}඀��PΪU7����QAe�e����J�֧Y�{�\��]�Z��	��Kr���lX�ϡ���G}�����Ӿ�h�?�PF�l��C�]�`Gm�!��=\�G�8������sϥ��h����~�%+�ddlq�$�^M�[Vwa�.�����b��KP�W��y��I��(@19�g�����7�V��������_�k�I�+��f��;/b��}7��o��(8�ѱK�����TQ�ظ�ht��hT����[V���HI����%�5�/1���l?G�i�N� �J`����vXR���o6�=T�W/��T$����u�|�GN�����:7�7ݗ�n�V�n�<�"55[�p��fJ�E߂?y�8C��d��>�:�޵I} H�k�>P�����,;��I9��������7�!<��t���T�B��jk�r!�ա&�,����ս�4�g�~�`4�f.D�
�`�G��\�PN�z1�1S0�||�zœ����h�0JI~�>d���,��m�{v�?tg�n76H~{+k����f���ݭ�0z@q	���P�I��0Xs!��ƳI:{8(�[��
��]�MZ���@�͖i�zE�æ����,�1i(q�@'�0��'CI2�~;��n��g�
ˆ��|��+"�ԍ�®�i�jR��rW3b�?9�+T��t��I��!Lu8N�z��.ض�,ͺh'���L�w��]Q�y Y'L*T�'iΰ���3��l�;陬	�=4u���a?IEb��=��TR~����O���&
AM�"�	��F���}Lnjap8�]��l/. Br����q|�;�`��E�͸�&@�mU����?���]�5�'b��B�h�Ld��s�4���}��"��QZ�L6���=h��kcs���J:X��E�-�u�ku@@�@I�&�0��a��	(��L!Cǿ7�N�fha�Լ��	j�h�HJ�K[���{��!��jl�e���d����<�H������S�G}k��P��ݔ�d��*�1ݷRG�����+A����~_0�|MQ��=�5Ӓ�)�<��3�%~�|���U�_��J>X�H�ݕ6��{�At�������7���@;X�S� �
p��=��ۅ�K��3 j�|s�/~�G��4�\���9�_M&���#-���t��X�z��'��&�wE�����yi�J�h_�aי�^O+M�r9�� �mx��PT��w#�ɖ�o1�k��?���B�� ��S�X@S�GP� ���6v_�΁�!���G#;��n�}�
��q�ޒ_:�D	���&�N���w�@�QK��h��_ϣz�`�O.�S�#D�f�/��
��7P�oU<��b�!�g���㰋Qr����3!��@Y�'(r�Kc�C��`���`����U�.�[��V_͒%$��*�������MZ�dMms�l��i"��=�IE�uby�)�58�x>q��%��.)��g@�s��b/g@1��搤$�a�/�����x�t�v=`j���0	�J��%�\�,z�	�d�[%��1����0���		{�/.���a��|ߛ�{v��s1���]X9~�矝Z��0;#�8n�7{��y�W��Y��o���9�f��Hо�k4���J�Hq�D�֌pE���=�N��F@�OΠD���ݾo�c�5K���v�g�`̲��p#|����,�<�ST�]�ђFJ<ĳCrc㑳h�����1ѿ��燢�=�ӔҔ��cH���tֹ�������w�� R�P����g�m�vp�Z�kV�&�&h�QS/ ���}^��PF�� �8W�Y�.Kȶ�<*����C�����0ԝ�����CL#���1�i�\��P�0��=��� ݧ�m"�ǏڌϪ:����4C�� �y����.J1:C˨������Ԓ��)�(��Q��L>���7��;uy���H�ӗ��V���2b�X�"�ˇm:�Z�d����Ҙl%�!�^�ng�q��@L�^�tB���I��J�U��۫Ne��갴�DH�����4�u2J�@��у�E�.�q>m�JW��~��g<�-#$�H� �)�i��NC2��<��D��أ�8�r
���q�}a��ʚ���� �2K!��i��"��Q�dۻ��@H��"���u�����9 �C��Ɨ�T�f:ڠ|�[y�ƶ��/�#)@����B��1�"c�H$7�nT��9�gӓ0x>h�\�_,`[̴ݗ�w��#�o�c�[\�Rő��e����^m�����+=&JK���Ԥ7bV���a�{�����T���Nh@v���@��PG�Y#O����矢�͌��Z,��]ob�b2�B���!��;��{̵ڠ�-[6t_�2�J�A�;"c��3�":�+��B�ׁ���+� �C�!zߦ�js6_夸����P�l�	v�J���hS��n~emn�I��`�x*�'L{Hvq�H/�^�f�`(�2o,�c�q7_|���76M�="�����:�Ǣ��L�(�wINlMך���^	%�id�i������c�,���j��#a@Mf�{����|+X����q��a~� d�����_}3�m(쁕��[������|���a�P�]��+|q~B������ջ��#����������*r/M�/���U���������IFF��3m��{���# T��Ǟ'�S
�/�z�7�b��ˣ
�������%�	���*5��߅������W-�PF�����,u,�e�8��`�P8���?Iy&dk���6uߚ��_�Id���?Sy�;�EWAR�
m�8��v�Ůp�h�&�N��y���YM�wQ��h.G��BZ�u���YB�B�V�B"r���L{�9�i�%����w�y�@x9�%%#c���>���慺� ߹��N�q�$KB=ʇ��WK�"L�����������7x����膎��g�KPR�a���o�����so�5dcKXu��S��/��U�VNh��_�)��!�}�ɡ��՗sK!�.Dq�;�a�aOc0�w�����Ń�צ��Gb,3�w�,�8����셑��C�Zb������S�2�xn��Z��`Ѐ�L���4���L����"�M&t�C�,�5�5�2��B��Al�
�!�*���B�%��4��o6��O QX��Z�T\%�5^�.w~���MjZ�w�/�����SL3k�3�������Z���.y���y���Q����U��Q�p"&��L|~/BzU�C�wG��Cpk������X-�Uڸq����P,ٴ�S�M�#7E���>�$�ס;���h&���T1�`^)����E'�ӹ��܌�f��̜��Ww��M�U��n�8�i]1Q���@jc�3�
�Z�3�D�ia���kkk��7!�f�[|!��������!r�R����؜m��x���d�1�T��M�8�H�r�s�O�9v�Ԣ���P��	�����"�~�4)�<�މT�������}�RO9	�7�+���6M|˼�wor���u��l�r�jV��v���cS�c�A�T3}�@�i��@~� �i�[��m��
�B�*:|��m'8���XD$�M���V@�z�7�0���_`�� ,Օ�A'������NP*3��@��;�CS9ɕ�K�T��b�P8�>����8Y{�CG�6V=��tk(*��sfS�c��<V��[��&���VH&���ߙ1)��Q��.�u�'Ϡ��Xѱ���5:�K�}m��_ш������ߒ��>_�m���QY>�^����c���)�O���?�'=��p�sT!�D�|���z��t�����!3��~B�C��Lo�If:�Ll[�*"�=��9L�6����k�0uz�F*g!�j��m���0o*5?�H<�ͺ�\���0�3P�6GD���D`�M9%2xH,I�S����qU~w���w�Z�1���(�+x�Qf58w738tq<�� 6c�Ks7lM����^�+��H��~6A����s�gH*�?�X�0���"$���.>5����CT"�+��e�P��B����ڿKj�3�"�<�FcNW�T��dB=3=�50��$�c}^��M�aM��L��@jm��kj?��Ƽ"L�S_��/��1�d��hn�|	���.$�T
��rq���k��vb,���Ŷi�E�x�g���z�U_l�ZT��|M�/�/���nx)�.��LG��B\��Q_�BT~�	J�pW�L�D�r�ߪ�Ժ~�;W/��&=eɤGz�ܮi0����Z��R���r�sR���s>�t�]I[9�/[LK�so���q���F�ʾ@�]?ZX$ݴ]�5@Qo������'���4ƈ���JWt�<b�/t���G��6�����&��}j�TBzڡ(V?}��Ks@�����%�Ա����}]���06�N�XG��$��\��Y23�8Я�'G�����*k@,�nxR��:�4��l�_@�`ޟؼq�|��ƪ���/N\>dYLh��YT���w�9~�ط�x����B�ϛ�q�/i����;M*փ$tˤ�J!����t�a��Bu�w(.R/F��s[�;..��p6�?���*
qq�Y^���?q4�@\�������Q�1K�����86Ig�E�L��V�o�Co�AU;��w�3�~¿aש�3R=�lD�2޹���(]Ol���`̺_���d��,�/�'�R���ɧΞ�WK�
��!kp�ʓ�qST��mq��8<�x�=%M�*� �U ^�Bw���/��郦�w?)�X�##�U�����273'Q6�|v˰�[��&|�;��Èޞ�ٵ�Ym}�a��Ъ$5�;�NV�=��cڜ�bi8|l�6\鏾l
��S����	���;nv��s�?�c��� �9'�]�3b�tL�]�F�zP	z��2�?�>��z��w#g��MprtB�ƾqi�߄����G��B[ 1'f2��;�9��d�y�f�2Χ �p_��T��Z��p�|ش�S���z=θ�"�����"�PC ��$�� �V����Y�������Fp܈NE�۾pW3��R�t���
�]#��N�;,��_������s�+5�[���z��Msy+,�M��21Gĕ�͐����"��j3����:�ɧ�;�ڌ�8q^�B�Η�Yʂ�v�w���Y�e}Bj���v={vo:���(I�69((��/��
��eavAv��k�����S�8w?B?����u��(뭦㏓�	*.^V=�U�u��̐�׿�2�^�5'l�
��:��h�o6������R��ǎ6��il�[�hϋ`so��&��K܅Y��������]<w�Up���g�-�-ސD�QbG���iu��Ȗ��� �0���&���\ $�S	o��;(������V��gA� 1��s�fn;Ĩ�?,�A�G�M�c&�8Q�u�Au��G�0?@�����/�V �'�೗N�!�7U���h16�:�\�2�%q�j��^�Mi'� S��t:��=�{�?�S	�=�u.&�t>#��`�@�z��cP5ٕ��M�O��990ݽ�v���Lph)Df�b���
2e}/�+�O	?ؙm'�V��8��6?�4�5������w��˚Oh�QW��Z��^���ӛa8Rr$�R*��qy��;)�x� ��:o��Vqa4��7� �����|N�l�wxjQ>�N;xI(�������(�H��,����Ư��^��'�ɳ��2?J���VL/��Jt��3Km\J�l�Xr��l����X�������z[�����*7nsv.7�K-d�)�r��i�+/3UJ�>D��l�a)�`�iըRz�*�Sv1r�ٲ��<�"4��a�0��xr /�����v�f���Rk̔t&a��/�-��K��h��5�a�>R�Ϗ������l1s��v���0�xuoNB�w�~�۷��t4&0E>�F�}Z��'�#.T�q��d��'pW��T��W�͚���AMt�|^:8́;J%�-z��
!Ƒ�]���-�d�>���#��c�* �����%lE� �1�]<�PVQ��Z����|�m���{_��(H������t�Z�D�x�VZ��}3��?��%���DB~`�	䞼�/%P��&�M��R(����i2�ʡn��⥋�u_Atl3�W6�(�8�u0��b�<�xb��b	�A]���/�_g�B��m�^�r�~����}U��7rj3����2)V&D����(��UbQ�e�Bf�� ���0ٻ_ғ������7f�m�Y��)�V�$�8"هV��ի�������[����U�/�5�0�@ɯ�~���8ɹ$N<LV¡P[?��n�$����v}G�
��NY�����Kr�2�h�� �A~�c���JE-U��}��{�Yq�6�aƩVR�}��_���H��x]f/to���"�i��m5��$�����*	��@�04�Z�j^L,k@�f�QӖ`gT�b�Z	�^��)MHz
}�a_��o��=|Tb '_%L&���С��b���S�r�6�^����`��@g���
;-��z7iR�<ڞc����.Klp"�|���p������8x7k��*٪���_ǔD?q�x.jn��[O�eܐ\��``l���s겳��ψ����Ud�m�B��^��]��}b�d��;*�X��b�ЙA` NVG��ѿ�'9�;�_1��XH:�dR�Z��sⱠ�8��:��p�->���r7/^C�R�����;6��3rYW���:r�{�%$�d9~��i"�h�]�L�;0=�܁G~	�� �d$���:6V��
�e�����y��#/��0wa����F��%���iJJ�X3G�n��V,�|�v��Y�PWs�[�m��=_�?��>��GFw��ކ����8�{^~��6�x���BD���U�~��[G�N���X�D�N>"���bG>
U�U��P�g��D��[0�Z|9莶�O��1&��V~ݪ8*��L��(��N폦u@����B��DX'!b�B�{_/���_��h G��d��ۚ� �Ҹ+~��M��em����Q|��b<E�}��O&5��o�ZJ��"xKx�T9��Rsxݳ�3�#�BClt�S�?��h��K4NE!�뀯8�=��_�6/~���X}ǒc�e����N�!��
���a������}Y4�Nͥ�g�l�c%-���o�?�S�θ�췵00K�@Nu*!�|��:�����*�UI�;&�By��R�,$Lr1
/���+J��b;�RźD�D�%�N����RԱRi�
����k��sqn��"�Oܷ_~]�%xGs�Q��Z%�B���P��<�{�^����`o�Q�=�^��ZpӁ���
j	F߃L�^bk���R��x�A2�"vU6�Gkpۏ�h��]N�s����
��?�\�}gD�}"ѬqH�%�yl KX&�}f��/|�^��q�S��Ol�^�奉����͠���	+<�~%��N���n2׶vUX&���W0a��ٛֆC0Y�oxF��`T�ƕSb�;�lTLy�����6w?p�v�+3Zv?��Ȼ������'��PjAM�]��M���g�5ˋlL�����:�~��S��<��Ϟ�[��.@a�h/���R'f�7�`绿�A���z�*�w҈Sa+�g���s�G��p�t�������[�+́�=����Y�l�[�.�����d�����hy�i�&Oyg+!$,Y�B:���Q �q'!���J8�Y@�	�ٷN�;	�>��8�&5C��%�`^� ����d�3�祤Uݵ����I�%�U��7��j ����>�``l����\ ��uE1q�
}d�����̈́�E�Y���H���:)n9�����J	N.������3�jB
���ɥGG3��G:��������
%Üq��><�>Z������ٯ�����k�&�M�XN�MN1ݝ<LҠM? ���6ų�!�@?�։=:?�hO�d��@����:͡e�u�����!��R2�"�6��4)�u��ι��.3<	�|L��4��1��y	��ጜzP��9P�؈����O��^i��$qH���=�~p��ۓ�C��B���1e�@	pGa�[?)q�K�C/�Uq�9yAӈ��j�y�՝���x�=%92�/'P���ɳH�H��Z�����M�D� h�
�|�Y�{u[kM��or5[��鋸
����\�4	p���n�w��Ģ[h�X)�Km%��ZU���"v1�d����A!N�HI�<�>�. T;�w����Qq�5�dPg�w0�<�9x�	�~94����;�s۶Jw�_nJY�ơ �;a��6��5xiH��R_� �~.�B1*�]r�E�gVm(,���:�_�D�$hʅ7b�u��q��Ή�m�����櫋d70�]�zmWz�`7��ӦN<D�rvu`�h)ʐ&s!�}]+��0�\I<TJ3ј�R�>G����F�٫��6�Q7�������:h@!잧������?�r�	2W����Վr	��\��:�%��KW>�E��>'���&x5��'�W=��h�v��Dһ�<��W��|~�C�5�3rz�7�T�H���|T��ŝ���9��$.^Y��ˍx[wh'��.K1�;=�]�y���[�+�O97�D@@/� �� ӡ~+����*G���$u�1yf��h��H��p�E',`�䭤�W��1�m��&����%F�-o^8�'���;y�]N�)��-~�Z��5"�^p�bH���(>Ro/���!�\��s����F�8�S�A4�	`+�]7��z��)u\�_��T�x�p����mb0[��������<ȖZ�K�'D)0;4%�P�$�wle�(���\��~Q�<��e�
JɄ�JP�=��p�@�]Di[̛c��}Оq��N"d&%��E,����緉Q8} �=�(��S��_Z����k�_���؇/*�,���⊠���mU%~d��(�pn�l�Zs�8T�s�D������ m�O4	��'�����|A�K;U²O���_�8�8Rrz�P�<c2]����f�T���:�%�FQ���av��3v���{�+lK�S��^����Eu4?��WR�GM�0�'���a��mv��%��vŴ�K,uk/��^^��ߖ������������o�~z��[�g���|{�o����Mt'V���?�������M����F��Ew!�F�Ӑ�y;�X���i`q	׳�7�imD�Q��r��*�I�Q�b�2��ɺ�erd�f�P%���
4W����hʬ���Ho�!{��M#D���R����]�¬�(�U�Zd���Ѣ��?�|]�(Xl�_-�f��2+̮�̧�V$�='�⦹��P��CU�����U�a�4�x�,�M��e�}PU���d���	�O����2����f�^���eW#0��[Xƍ�S/��,g�F�V����orD.�ND狗+�8&3l���3�#T�ad�Iq�~���W����_��p�3������Jz�AG�B�v�������H]����%-�f0-�3mO�+���m3伶�h6��>y>�7#XJ�*w�i(����.��1
�$�߷�2B��LMF���4TƁkHw' T<'+���m��_<x(�JQ�:[u�M{��HdBD�Z?$�lz���`R���o3�ۃ/�.���t.a��'����Ҳ3�H
K�QJ���+�4�)4Lbl#ܼ�ė�K��r���g�
wΪ�T��J��r�β��n�Eu��Ga_���W��#�()B��K�@"���j*�[|�Z�Eg03DȢ:�x8r����T�톽��N��;�zl�x�˚M���&� ��D�݉�J��+&���F�j�6(�-��e�r2�K�Wv���zLw�@��6�a��A�d&�wY��[Z�)�`�M*+��mS�p"�h�K������h���F〱-'o"6�-)	`,}�0�@�QO�#Pr�	t2���rӟ�W�;0vE����%��"�nmԤe�E�s�;��|֬�|�]����S;f}�R�(�{4A8Zq��Ӧ� 8H�rf�x�����]�M�����v|��m��i7���9��ѴXN+dCP�e�JmI2���$�;�p�7�>�+L�� "5�vP��@�"u�X1C��Vm�KwP�9��ک��d	�ʾ(�9�m�E�?PQ�`����r���4n�2��?p�������/�v1����تMo5Q�08�SXy�hXoZ1:���7 �S>+���2��f�+
ˤ��yV\Z�u��Y��.�p�x�PWr'v�G�.E)��v�GGtl�7K�$~B��9	��l�>��h�;j㳁�}R��9$�n{KJ����\����S���2�у���/XucZ�:��狹B�jx�;=�86��<���M��5�ZZ��L���x��,?�Ptf�����tReô�Q�NQ`2S���?�`�Ej�O����Ht;���&�)ߣ�b�#��W�5�OB�euI�}��.@���1�/���8O0As �Td�/�v����wem|*�-���TJr�������:�C8笇��h"j�7������w1�f' D?�{G�xll��|^��\�%{���PO5����y
��TB�l;a>̖����D9��i֗�h~scצ��WV���F��7j&Q�O�d�iE�U_��+-g��xw-n�s���7#1�l����/;�q�$J�X�����T5���Ľ�)�� ��� ~�G��l�;ù��:o6�����@���KF-�^��K�4|��E�	]�3����FŘ|A��id��s��ZNw���⭘�љ�o������8�Ǩ��A��_`�:�B�,M��F�3T/4�������+(���_.&��x|eRUH�O*�2�3�u���Q­���s���#L���`O4�7pW>�D�o&���4ΐ�-<�U�?G3��j�8Y��*�[ͨ�J�����w�:j�6�vƳ�é���6�+����ԟ&R͢W�l�䰓90�e5hlCSU/4CV��#vv~���]6��]%,h�f��]x�Ŷ ��	߅q�\���j΅�nKN�G\�!j}5ϡ�S��oY�t6YG�U;r#�� �<�g���A
�}@<�ߩ.�fR��7ʺ�8|�dùE�o �-[�!I|�WN=C��ݐ0�4�ë����
9┭��u�U%[5�w�/��(\���$���@U'S���s����� ��Ts}\���r�v���].eZ{/����ݮ �a��#���m�[���"����{�S~�bNW�v�>��!����rɖ�Ɔl�5�bx#�����0)^���mw�O}�G$hhC@Bjn�TM��za�<��Å�èk
*f)Z�x7$g�+��$��=N�F�Hǂ� ��9v[u�����U��S�2���u��j]��F�fm��,[��ɣ�2�~^�o�3z!n\yS��Al1ޫ�	�;���3u���%�Y5�~TLgB$���sjA��2S�p<�C����i����֭�[�S��LfVv|lV�47\��挖I�MSx�0G�ӹ��?��W�eġ�˃y�!�OF��6���όx]R���l��i�O���4����D�S�~� N����w.��*{q�݊��14-P��4���u�F�w��]������@ιb�j��@BN�c�Qk��NYQW�qGBB�\����OJK7���@��\u�Sٱ/K���Ȧ�ۥ������N��DD��l�����fj���-!=�¢J�w�Q�|�:c�u�������ƺ�\�3�4<�i�[j0,I~����@��x��˱���Ya(��o�*hu?�39���UЕbn�������:��`8JI0��d*��&���b���c�R��ٸF���b"rp���?���Hҋje䘠�����u�?d��G����U ��L��e�_!k[�6�Z��"��a6^RK��˒��P�g�֝~�4u�}J�����͡�i����1��z3=����������n��$�6���M+C����m�G�JmQbk:�`��E �?a�`�;��E��<}'�@�͓(�2�3��D�|2�)1,�^�P�ǵEeBm��mp����l�����9��4�1M�nè�/��p��,}����~��]���J�����_Z'?�z�ި<���2��r!�F�O5�r��e��_E	� �~�vA��m�:a��&���^��凹kߔ��`�s7O}�����|F]Ҩ|�16+O���H�!`t0�f�8����͇p�ɍ��}7�]�]�����&�vн{�\��V8n�����̍��B$3l"��n����������Ǫ��a����jۿގ���ӫ�˼1�8����%��hC3�ʞ���Ǩ�{�.O����T
�m�.f��	T��]z�Ư�f?��}qs��� �n���:�]��fW��b��u��o�\sn�~�������C�7?���7tP�Ok���E�_w����*S�����6x}��_�:���b���k^W�oN�����!+{`��!�`�=�e��}��7�CAhh��y.�^@����B���:Z��3vS��T���>7a5	i1��r�}��Oթ��D	=*]��{|�q]P��s�'����@^��9�F�~t�xTӚ�� V}F������e�C�����z0).�;`	��_p$����^M�6�|�@jNg�"o�������\�0�>�n��.،_�Qtx:R��N�ּޯj4�� Hu���^���I{���u��^i�Yk��7_C�iE�`m+�8��;>�!Q����,�9�[��o�]���j�!{�
E(�]�\�F�v��#�A,�Z%;�J��G��!��@-�H+�Y��5�!��`��[)ǫZ�qd4��GZ5l5�^��@6 A t1e���so�'�Y���L�p�_�������Ο<����}�	��v�nq��d.���J���lz~0�oӳ1�4<�uAծjx��Ԇ��������W�p������=.�Q�*�>6�:����L�]�ۚ����mt����*��?�1�tw�<$���Xk����JJ�*׿����ѫ�=AF`�X���5Fʭu@�E�yY�l`��䳪�b��cslY���P����d��^�C�\eED�{��6P�]������`���\�yA�|�-���y�r��yF��Mu�?̽�I �4�*'�y��������c �Gކ(\5j�8�p��ӕ���h��1F�)�Jc�/�C׶����=ho�K0�뷱�"�y؏�nߩ5�%~�b��Z-��%�6\��y������L��긖��x1�?�鉿�8�G<(`j��&nV�;����b���b��s�j�\�`���ٙ���y����F��HG1�g*K��������o��?�Axb̜�#��M�'�)��4-őR��2WGdP�x��#.�t�G "��au���VX�t����<�)}ѽ_�kAv�����h�FO�;�;�f��G�w�
����J�Ji�7	ח�o������b𰢔�R@��BJ��dh�]�o7��)�O���� �|S����;y=�43i
`!���1*���M�%>�&m�Af�'` ��+��D�>��H�ߟ}�Y�-IO��!�U+���c���zj`%�d�=�x�jPZs+�) $�4����n<aEMUS$c�y�o�������j_��UW#���2����8)P�H����ي��3�N��E[%M��z�nXa�S����;p�����Z��$c��V�O���>Rq��Kg�:~�������O��!w�"	.���K��u��+eүs���2^�@��6u�e�ĳ���kw���V���¥�'s&�{9�2��%Hט��Qx}�7�[0���
��MЯ� ����\�� R5��^��0����ؖ$�70����R8�H���aB���ˁ�����НK���"Ws����͌�_������[�Jze'�ݬM��}������$4!�Q��l5�t�~P��B>�d�8yl�e��V�+�$-������,]XJ����c�z�t�{wĵM�|�e��¤P���\���{Zc�o�%�(=T6=�B��8�G�E���mT��671C��Mℶ&܂�"���+0�>�5!e�H%������3峤�B-=�A�%`�s�r���/�H ��]������/�˖��f��a�j ���Z��+���b7%	����e1HS ,�(b��'Դ�	E�|�=4#6���rL��i��;o�������(`�4(�t#J�t7HHÐ

J7�����twI�"%9����}�����<�޳�^�z�s�	M۸ y���=$16=~�MD׹�Y��]\�������S���j����zO־&��������f,���knvT��S^xX@Oz���#
�8*?coɘ�(/�0;n��6�W�τ���v�`�Ӈ %��.!��(Z�5	U|���;�Ʃ�٘Fމ����8��O�od�[�)�}�s7�o��Xº��g���[V���wp�0��$�����ǺQX�ndf����'�뎖D�8���K������?�l|y��dV�-��9����g%��>:6��W]��E��M�ǋ��b�O�>}���t�����Z�-�@�U7Ǔ�s������?�/�/�H ^����Wy�qj�|a9�Ymi.�:F�����7�9�Q�^[ο�����*���~�,�S�O�cϷ^E�~�j8�S&�ix,I��E�DR6F����{R=*t_'�q�Y����@�n�V��I!���5|��ծ�X��RT��o��t���K=K�"n5Y�V�72vC�?��Me��D�\�lsS�͠����굄67�|����|��}�b�n�����aVo?}%��c&�Ocu�?��U�ң�p�;qͮZq1��Y[�HJ���w�����p�JZ9
���@��:uy��K�Ew�Lc�͎ֈ�
{kRa?�W����)��}]&Yx.T�����MjU��VE}}7u�n^��9�!�]�dhw@r�(u�q����3������l)�y*Ns��Z��&�7oD�k.��W=-UϤ����괚�uܔ@�`�-fxײ����&�S�*P���)$���z�]t� :�IF��W���s��Ȗ�6��V3��G/�h�t�y���J�_�
�8�@��d����������Ld��՗̸�n��+�CN5>��K�D>�1�������F�V�Ov��{�9�ƒ����$J�^�h$Ǹc�i+W��{�iB���u��Y��g*8�St�,Us�y)���m��4�c	���ӄ?�<J���_`Pz���ޟ��y���t(�-�=�˦5��p�ha
�U��3�����B���z�j�A�
ߎ��g^9�qCOf!LM}������Y����t�M��#C'�|�߸T^:�F,�3H:
����C,q<xL����y<DRۑ����$>{mHyܓ;��>D�y}r�=c�B��߿k�bF�:b0:����v��;��!Dd�_�3�<��|ˤ�T7�ζ�#~OI����><3y�\��O��~��-�tu��oؘ���7�̱̇v46�87{����~.d����]:�:6��◑����M�Ԇυ[�v�����*����2� �	�-����](Ƃ�ݹ�sڵ>���ޅy<���j9ӟ���&3v���H�)W�c��;j���k��[�x���`��7?c�`��>�����x�~�祪<��?��[��%�/�bz(������wދ#*����7���>���"y�ƫ�hTqM	�dx������j��$�dz��Ø�U�7/�=~��A\T�§������؟4	��I���&!��<6:
ݖ���1o��ߒ��Z��R���,�k��'D��`�t5>���;�c��:4�S0�>���?�'<�����F%&���c�+��Z�11��\�SX8�ӌ��}����͵�ۿ��|��M��}n��1M��H����[Ax�S���Z�.ZVN�YA�G�/y�1}uKu�'�n�=�LQ߆�E|qƉ��	N��PJ��e� y��=G��H]X:������6!�<�_���XaD]�8�i0��tr�l�թ�E��6���0�uU;��V�xU��'H���*�yu�rM�^�<��/�+_�U��;�lN�_T�J"MjC[�O�|h��V��V�uj�rde��[�UL�[Sk���	Y�2(�����SM"RA/m�#C�յ���ߏ���{1ʨ�R.%D��򨱨��O��xt|o=�+�Jɬ�wg���%ɖ�S���6�ʼ��[�+]�r[8�&��O���V1���Vʱ�D������Nq���*W��f{�z���z�y�A����A}2ns�3kYPGN�0�궜�Mmf;��*X��2+�#M�*f��Zg�X�o�0D
ON�c��5�f��ڇ?r��E	�b��k�>�cƽ�Űᓢ\�� -��Z�˂i��N������?����C*�u{r^��p�mw��;z�x�7X�>3�:���f�4��@d~����B]!�q�̷�)��
���Yo
#Xb��p[z�(dW�r'tn��oจ�бo]��x�۹�����},bJy��[߀�nhW����w.��cQz���|��Hc\�H��9%;���K��Ym�<Y�o׫��,@:��c9ť8^���<eT3T�~��kf�zm��,1`~��qۤ����I9�σ��*\��;�7O��V-�/��/�?x��2ʜ��_�b�?�����@<�U)ӽ��<YM���.��t�rk���3�O��q���`>�\r.96r�i��蘿24^S&7T.���XIt����Z��b�V������>��v>M��,�^�M/!*�'̖}�m�0_bM���YNG)~���Dc⇊�5����&J2�)�o�bN�{5�����I��_��9�?j���v��N �ش?�����$<e8@w���X������"�b�De��2H�9���b]��l��wF�[�A�"A�3.����F�C������W�/���&���M��c�����Q���tc2+ޘ��VHv�]�O8��]t�^���DR1w*��w�7��:+��Z���V��կ�;^[X��Z$X��Zl.����a��
���~gw��t&��M�~II9V�X���@O��#�
���}G������ˣ$�9������������To�>f��̧F#[c�~�"Ĝ�$.:E���F��x+�kSdh�?�FS��u���,�S�YՑ�G�Q��n�5���R��ݭ��fUcX^��|��w������cJ�࠶�=���t����.5N����JPQ4^�e�sȹZ��G3�)#U.ڑj�2"��l�,���ʱ�y-J�	6n�T��.��m��B�r����������v¬<���%�S�O�̱>�Wc���AE�wu��
Ε���Vy���o�ꝕRC�tcm��~����4����7#��88Ոn��JĠV}�p��
U0;�`}~�ũ��Q/f�d��01kc��G΂l��I&�b�{2��n[s����RS�����ɢ����<����B�_DwĐ��R;( )(�u�>�=i�N�4��O�x�2zu�d"+��b?�J�I��AlJR�A�t�2�>n}�LC��=�cU��h���$�De#���X\�p�P��M=���K��YZ��5��H���1:5��xd��2V_�m3mܶ�����:#�����.z�ZЏ�p�w��C��j��Xa�)�ʙN�fN�x��`�\]@�"�&�?챯���%1U��|D�EC[ڷ5"���<���ny��ȃ�==�H��ȣ��Ѩ%k4|�<��<�=��p�]��}��d.81���f͝���$���ܽ�i�U�a���t�[���F�9A�`���i���'�bv����m�!�7��p���{�덥��͹��,��8��8��sZڠ�?a�{�/�̌�Q�cQ�_�U�]��3��=s��ގ���6��%;�2��u�E�\�!��>�� ���Hht���F�Ռ��$�LD�:��?p��DF���ޛ�ټ��u��Qo��A5	�����݄GF2�����m��~���>�h�9mu����}q�i<u>���np·N�~��݋<O�H���v�v���Ѥu���.*So���q���پ&\��bT�r�&¶�(��u��[^>�D�t��	*-��]���9fl]�������������? m�T�v��M�sE�5�W��ۃ/U���3��ڧ<{y��Sf�3nPgUk;U���S���/�'<���?#N�p���w�m�ot�i���d��ݿ��|��㓆��{.nl�(���]�w)�Ջ�
�O�Rɔk F�%F)��8��s{�R�pI&�V�����y�7?�s�S� ���&�X����$�Hħ��ãN�;�y0��Ρ-��?�M���o&+~3S.�3�0��EX�70)>���Ly!$�천�O��i�Jt���<+��%��Ʃ0���$s��9	���`'C��q!�~�O;oE<����vև��B���U�\@�q&�jk�_X����5Xl�����|���,B 5�Nc�9nj�S� ��Ñ�r���fM��	���S��W\�P	�X��V"�v��7A+&:vc۽�{��g���uR���E�Kj< ��	֎�W�?��)�.t����o߂!�fE>Nm���'�K�����b��Ԯ}�^�R9�d�������Y�2��L=d���	C�I��l�AWO	��<���0�1�S{�������-�ӝr;I�$�!���p$i���y%4�,,����f���h��������a�Ɠy����Ӭ�d��`�Eo~���<ߟ�v�k?����Ie�\�;�i�l̞>e/e�̬!;���'U�T�SZE�OQ��E�'$�j���B�˟&Mn��0%G��w3W
�p��_M䈿�� �2�{�i�x��XI�WݤL�7�jؼ�xґ�%�	�V4�/��e�+%.���X|�(�#10vprZx�7?�'��6!!}W�l昉gG8M7�sҧ}��Y���%�R^�L���ۘmMs��e����ԾW��I5V��+������e�&�=�����Ц˟r������D^T���TGl�y���zk=���G?��p.��/�Bۼ�j�'�D�|�9�(M�w�����}��5�1͝ʪ��n\F'���=��=Sw����v��v�د]6�oy_�e�\��i����dWgd�L�C��u�wzZ!�'871�.����ӏc��%�jx�	��0���E6���*7�ׄ�*���'�*���YC�/�x8��~����/����53��(�Z��|P�M;U�uڦ��F'5��}��e�T���=��{�m��U�
��:/��	k����t��Wf����*�*�n��jze��I��佃��ťÏ���.�
h/�tf�LŹ�mf]�����B.-�@%6�7M�󤀜�Հk��ҩ��W���@���
0��ݴA"�z�6C���>��xW��0?}�$�}��ϛ�m�-N�	�(#x����a}6G(|�骓����ˤ&h�k8.�Ą�ݖ��l����ёYe�Uf�H;�����q����`�[ǊvJ�-:q�u0A�����^���cs3���~em	'e���i1l�G~8�9I�3�|�8�����s�f&���va#�/b�7�k�� !���{[=�(%1;;�磬� ��pT�1q�>���������@q.*Ӵ�ʣ�XS�l<�K�
����k���?�?v,e\Č/�J��������$��c�6g���&ҋu��7HxX���=鼾�|\b�<�KK�!��ǫ�(�1^����b��1LQ�Wg�xNwwu'e��ɼ���xp�|�=�����G��IV<���Cީ���+;�W�	��F�aL�U�����!�U��i�%��3��V����-�#��6~*��)�ͤ<�
-b�u�*a���mlb�nP�IE��z��H��,����4m�d����1����|+����a�G��������1�n�Z.��*y�%��Lԣ��K��Se(�P2�e�V�򠭦�]�)�����vx�w����lŐ�77mm5!O��G��k�R*��8mV�o��:��Z�Ʒ��&�,3����͏V�b�5�������Q�������Y��:����bu�����j#������H�a�����'N�o��|�qRT\�������M�m�(6��{mq�Q���+&��P��ׅ�#�
�ܸB�>��^�QD�ʯI)���`����}��{2����@	��.+;�lb���8M�R��C|yKZ�@��;�'��D��!A*hNi�m5�1.�e����D�T�u3�% �4 +AmKo>\T��mt��������?8�Q�ܭ����m��L�9���q|��`��������Q��r*�n1�{3^�L��Q�z�{}=�a����OV�[�!�^���@!r�Gf���$s��j^N�ջ,���e���OiB�x!�7��aU#�����r{�N�f��4εk
�R��*_��.�F�������q�VF��>�ݠ�7'+����;�ʙp,C+�S�!������p����|b*J����Q@���py�y3��U�r����o�a~�Y��C��G�pUk�JFH�V�{�4Ω���`
}������Ӟ��m�.3����������������E��tGT��b���c�	�F��o��b~m��3?���!N@�fl�z'���ډ(G�j�=C�9"�|B��q��?,�[/�zޤ!xA-��l�]��sX��K��i�hH�$uy
>%j�����'�^5�{o�,�Cb\C*�-��^�Q�aV��l�a���b��:����ޤ��q��:�2$G�Έf�|��?�U������d��&ۤ�S�;��w )��?���>G��s���7q,[���fēS't�����_=Q�#P��T�H��/XR�U�P"P��)��pn� ��7�.��\���5�ȹy�����Tp����5�E��qԛi5=c�m�b��T;|y�����suv5��v���'9�߫�)�)~�6��Lw���]R��omJh8��><I�,:j�4�=�dh�A�\�ݡ���g�~�]e��2�S���ÑA}�>,�vMv�H��
��(�sd�>��{��;��q~��l�f�W"��;�j�Dc���"3�/<6Y�w�)��ww{i�T<���_�L�\�~؀�o�^�B�1UcMv�N*�B�ٷ�t�2�+�a�
���"�u%1��U�89�{�����:-_�R�W��֭f�<��lU�8��"�6Ȼ��a~"�a�1�\�G��z "RY�Q����W��&���/���6�r���<�����$fH|�"4p��1���E�<���c{�q���˩��F�{7>U����w~}WSR;�S��vm�%#������<D2�N�c��S)+�0t�<�h��÷��t��ԠGx+���qa���44����B�X�:i�j�Χ��]��c�B��G7?�]��-�V���}�ʓ���I�	��1�����B?&۰�4�I�q�Po�6�:��٬���܃�I���/^D� ���dv�ګ�ȳ�uk�yI|Uq�35w؊�̌����[rF<�֡ǝ3V�s����>rrP���
N�#�2�uC������/>��O
��+��?5�7O�k:V*(�	]!wxp���~����"�6�lY�������`մ;^12��]�l<ˣ��(�Q�n�p��#������$Y�=,w���gj�^Z�9�kq�8c���0'5��cFg>���~|�\A�/Fه�CW��X��h}�̀�"8� ��:�O��ޘ��5�q;S����2�@g�9���oZ�����?���ˠƈ/eT�#�F��Ј�2/�[�4z'O�gZN�>��z�|v��w��y����D��҉xn-��5rf�f��#O��gc$"�q4�Y�i..{��zm��E�x�:ǥ$�+���]��!7����yq&(�Ԗ���S�Q'7�������*K����iFO�u�P���B}��}�w�Y��:E�?��7�z'�)1��&��{���p����Q-twůuz.�)ΰ�1�1�T	���k!���-M�	�6��tULh��H�7xT�%�1�j���x�Do~�YP��H�T��~|�r�n̬C�^�;�*gt���rZ�0�b3�������&�k�s'eU�{�54�{F\�Yq&}�����Ȼz5�*Ը�����mgt�ͧ�~��+���fB{S٘�h����{�T�`(!�#��a ��r�\_�b��Xsd�|�ag��ۑ2�VY0[���Y�z<UD��-5��[��U�j� �Ky��:�]
f�l���+�Mq�8��)�zK:r����?�O����wR9Bש^��}���l��)�Ã���P����|R�G��Km)E�4ך����ƥק���i�}��vW�-�=���"�>%��M��gC��������,���� $��pZ�KPA�9$M-'tV:T�#�>��ѝh!�(A?���Rx�}}|��'�B����)�:i�m��������2<���0��С�p�*煔��s�o�4��}Ǚ�+��q1��C:�g�)�o�]b:�*�\Jz���˿0��m�6Kbv'��b�F��;Ű����g����}Ey4ua�0�pY���ZԶ�ɛ;���Ib{�����ua)F�Y� �_9G��/����2H��C��ld���겉ͽ���2���5rN�L�QL�
��SL��j��y��5�y�V�s�+�����5-��8����?s��u�'�?�����X�J�S�NH;q��ؗ�t�{�Y���}�R_u?]�8᯷��$��K�]2�jB�`�U��+ .�wk,kvj�J�����i?@|EI5e�+?��Z4�ߟR�{�߸aFڿN���ڔ�����1?3$r�I���ה��]_����8Mv�,YN+��r���{��ɂã�EčYC�ۣ�.g��:�#��y��^���=��ܗ�Ñ���͈?�棯Te�dW��;�L�;�"�1�yL�'�_a��b��j�dN;��x�?,WN�]\�r�P���!ts��
��t�˭)�X�Y�'q���ً��e�+��n+g�z��(:�x�BT#x^�oc;��;wH��g�� }���Y���f<��~	�Ǆq�}��@��*��K���:;b�r�0�qq���Ͼ�S����>�sw�c��ɘS(<<��(E�����뽉�(����:���������~�k��K�OO��9�z�rJF�X	��������Ն��p��^����H袎��)��u/SK)�.�M�����*0+�t��"��,Mn��ɺC����WrΘ4�2����Y���:�U7I�2L�A�Q�a3��^���I_�mxʉ�KV	�� <r���ֶ�7f���4��B�3F�3�4�ē� �g�i�O38�D|#��	�V�6�>�����,<�$������ڿEJ�2��	2.��wgrhI���IQ�����Y_��cRE�L-)�mG�1�����6��m�/�����9��r7��z;�~�$���852^�Q�ԗ�����O^����-����ˌ���[h�� U��ZU�r��b�1��y��^��)��7$��~R���w{�GY}2_��~B�/8�4n,L�܎ߵ��4��u��a��8b(Qg?r�W�r�9����z�J%\��૮v���h��M�#���pz��E�9�6�J��N͠�8���,��:�ԕ�X
c"�0��B\V�4㆏�*y��^�5��N�_<�����:��څ�_(��ñ�"�K���'�z��g��Ky�BiEt{�����I��p��ҋק͔�	�'KbQ��/�]-F6t���jO�X���[��+�ũf>�&�G��ŔToB4OĴ+�f��ʒ�H���qDǙ�/��5�܌dw�:�M�:��*^-���1d�Nh���})�����y��t����Y�Gs�
a,d6#��_��-_X��Y<�{���sw>e[g��`S����%������������<r�P�2����C�}y:� �Y��*�]}�h�:�_�hT�i#p1�]�zw4��&m�7�������s
Tz�4�i��jǜa�`��bͪV�^V�Έ5Y}���:�b}?�a���.�yu��N�������%/�96)��)]ZШ\�&<�IЫU:���7���A�5=yS̧k����υ.��0+�j����f�ph�S.vcڇ
�t�D�+���N�o�l�ĺ�L>>��x��Y|��M�,��a�)�g���.�W-#��A܊��"���o\z�e��YO��;t�6�,�GFgyđ2���t�P�M����=��,j:1��{�LO���HZ��pqKȓ����4�=�����WF�ȆhJ9}�����9Ś���6�@�>�$���/�������0m���c�X����z�bA�|����#t��|�ĩ��kČWZWX��uA�'���ߓ��t�rs���g�>��]Я�cE�$�l8� LFW��_�NY��S����e�}�^e�=;�~����_ݼ�̫��8����t������F�:g<��.`��O�p����]��$N~�����ߡ�-��b��+��t������ڒ���e�UK{�Y���]s�g�����8���Й3<_��:l�xVYF�%��m�-tc�qŚ��9�I��.g^�ý�G�3e��"��P�*�&'�>��t�5�vίn��5���*nP-���ϼ���l6�^�� �E��E�v4�_N8�A�B�%�y"?�lը7kn�H͏�I'�6Fy�d��[?����c����K��(����=�U���c������5˧x#��I$���(Q�K�<���wl����ņ1�V�/cB����������n{	�B}�"�x��:���y����<�z�9�9�g֧�c����sT�I� �w')c�a-oe%�g��OF_�Zi|����gG��A|6���Æ�g����*s=x�2}[�	�{���E�|Uu�	����W�1�)c�9@=wb;�:ɭ ��Z/K���ǳ���D�#��r�N�����$�&��5�[������T���t�E��
#��9���b��#>�����q�>|B�)9�s��Y�5�!F���/V�U��~P8]�ిҩ
�]R �
a���z��W�L]���q���Rr0=����/�D�x�D~b�FS��	yK��m$�0��oؑp���ql's�(
�Z�6���k5�2�ۓ���/b��	<WR�P�oj,7���e�C�`��Ҙ*���,�� &'{����B����LYp�c��5rkh���_��0N4H��R%,��<z�EN�.�޶3ۯ�.�%e0��b&9.�8�d)���W�+�E��"���Xd��M��Ԉ� Y�g�Օ�\Q�C��MRv}��ի���>|J�[��es(I�ߵ�&_��+v��z�|�8��$$���m?ZkzR0����q�����T�-�uop�?�y6�4Qh%�� �yw��yI�>���a����t��ƀp�UH=7�P�a#?w�[Ӕ��y�̃GX|�sD�yʫ��)g";�Q�.�4�/5�w���)}�٬˥�Z�Q\Z8�ܨ�b�� (oH����oq�o׉J������e��?��8-T�>�S���P��n3k��H���͢�w�����j#6��?
��R�����<�9�'7uʽ����I��#S8��B�m���W�)Y��' <���������_^���l����B�G��|���F��o=�Mܪ���щ/LN��u���u����;��d�^���Xmm�z�;��^�t.�ը�m\:b4�r���z���޴�`��r��P��>w��ǡ�Ja�Ke$�pE��'�N�:}��"�]!{wQ���i��x3}	w+f���!��+C���T |B�7ڊq��I����K_�m�������y�ҁ���;�6jY.��C���i3���s�v&e��*�:��(�&�~�������R)N���rM�SX��:�~�'�qt�������Fc��5~��:�5_�������%����^<֯Ҹ;nW8�S+T�)�٬�?��y��q��g\Dw�#������;�b���]g���1s�̸GNgU��Ow�����>8��??sW�o�U��Y��d�J!�^��Y�O�?�b�4�g���6hls-��=}��Ӯ�?�̡򬞶�i������a'?=��|��@�~2Y���ϼA����O��tI�!�^+��soefn<�Y�����@��oV�bVIG3��w�V8�Y{Ud%
O�{�R7ҀX틴���m��$:�:#wx���4�i�Ġ%b�H[@�]���u�D�:�qjkp�hܸ9*�aщr�d�vtq( �w�R���X ���ɛ$�������.(m���B�:QQߴ��c}
:��o����k��s�1	��:ۃ��Gp�|���s�	ڭ_r�/
+����r
�V+��,�Q�mj�$�H�������W3�A���=�柃SI��'�uRw�mgS4j"E�8�9e!9,R#�'���������2ES/�T�%O����d�kz4BY��ri�aP��rpl&['qX�CW�K�����n[�|٭���=ʷ�˟��[��J�Y�l�'{�����6����ߡ
!V}Cr++����mBWt����J��#�2]6r;O;!G�(:EǛ��sOMM����b���5��g ���ܓ���fe��켘��'q�'��'�x�����5�;e�a3���ߋ����7�uI���ao[��Y�n�F�t=M���@^}���O_:QQlp@�s t;X��NЖt�����a ���ã�napsV��I����fł��+�fT�,�f�Px˒�#��)))�w&���@Gx��I��w�Z	�`�Fڒ�m�,0X.E�c��u�S7� b���:��yi��]Ip�}  ��Ȅ������#����\t�jb2��)�{�o��b*F ����+z�A
$D��db:�6�5%~�b��H��E<�?+D�EhI�PK���j��_���f�ڄ�m0XY1�>��k�7�u~��th0;��+�>�E�Y�<���� 
m]� �]�(���h���8�x����f�ԁ���]t� |iSh�'8������6"h�kPZ{�ԳX3���E��r���4+`uq�+���#hl�b<��5�i��GP7�n�o��]@��~�z�v�G��<�P�"'6y�9&����F� H?_���h�F ���`�⠇Qu)K ��Cv�
����J���*�����E�r��D����q��wP �_
��>t/�~�6�������z>��Xb��8x��Qy@ކ'B�3�{{E�D�A�gH��+h��dm�b���{9��=t�������2�r^l���5^:D߾
A!�=	����wB
��ǋ:L�3jї��z��C3((ͮ&f�6�� �H)����@��?��E�`�3�n4�@sL@���p�wL��4
�OB�Я��f���t���=�H�R0U�T��~!�G���)4��BHp5�r뷐��=� OBH~�P'������Ӳ�:Y���%(���@Pw|��4� �y�q��2	�,@J��0p�&��:�on��n��&�P��nyI2�%4D�D��`��A��Ac'h�K��F�Sh�$Wv�Cy��x��� �eL�� �����560P�!���"IVP�DZ�� ִ	^h6�-���!�w@�a�ڄ�Ҟ�(v��Ӣ*'|N݋Y�}"~���`� x�����x�Ā�*�֖~"������'Y�	 i2�^a���ꠜ4���6�������܇2��b
�R����: -�@9���,_8_h7H�?��,X
\c��H A�i����/A�^���m�א�p3�O�`�S	��fK0�EEm�#�����|��	���Y�O}k$�
v� *�*�7z�� �O��s^�r�훐D@��(���"�w�+�?�e���!Y%�6��i?�y��t����C�x�@�
��W�Et���@���!�	y���~��M�ߓ@��O���$=U��%շ$  �x�� P\7 a>��A��0��m�.�v �)��4{=��!��>W,{��6t2=��)�����Ø�����i�v@�P��ڵ'0�A{åe�A��~�*f�� �y��4���K��^Q�2�xC�M�@�������& �k�
��.� !��������?	]�xE!�ݡ]:�D
,��ܐ�w@rCDJJ��r�Ȳ	!�����@A�M�[' B��f+u�d0c3mB0?�^�8&/�H � �!�/�ԥ&B؃�:��8 �� ��%�X	�n� ��� P��ă�eL��ǐ�!�9@�(_�%�A��.)"BA��Ϟ`����	�/��&��, ��P�@����߃X|�����A���%ȋ��7c_y
p��+D� cȪ�mD����
����Â=ć�����4���C�S��j����0��20o=�|I�:q�P���2�?�&�!�K���C^@O�7��#�q��Z_͘L@������Rt�)���w�S!]gC���Ѿ�?��q��x�y-<����A����}������?���9{g��.ĕ	�z��N�$��! �2���{���O(���/QA��k~����7��,��ѐ ��x��J!k-~2�tl�ԃ�)D�� Fӂj�Ex���|' ���D�פ���m���4���q�W��xW�*��W�3У�����������m�s��B<�����FA�u�Ĕ ���֞
��W"�5�{xv������;Z^��$!�����**Am9A��֒�P���R�?kWu��讦�Ax�0�	��6ӿ�v��?B�����o�-����?k�� Y	A�F"��������]���j��7�i WX��'�/L�7�p ��m)�r���C7)��:���hf�\'W���2�7o(P&ea����i8�n�� �P�U��(5��ǂ�C��v�H$���AEf��MЍ�[Z�G��U|�� ��[����qKY0Y�'{`B㗼�Y�gP��_@��������	B��
�%�q��,3�L� =8/_y�U��R� �<C݀��~"*4Q�ԃ�0*77�|.6��@�����io�L[ �	Hwm}v�.E�&�h;�A�%M�r�	hI���������#ٟC|٠���bA�_��}�"�
�#��
���#"#-��a��W{'A���@�s;m<0ڪ�e*�d~*G2�*��|��Dx��ҭ�/���C��L����N�F�9\pa����m>�����vl�O���-�t����ꂜ�5К�Z�|u�ُg�6!k#6����0ns�@"����tV�jw �\U@؏_e�zq��|�j�����5)U�KѹN�a�EK{�^�oHF��`���&/��o���o@�ܘ��X��_=@x��N� 2Q [7�J����9|�!�	���1Q�aO�^tM�:��w�l�i�[��c{�*yi���Y ��L����Ś���	�l�����s��8�8_ FC�.C��A��7�	x�խԗ�|:�LC4ׯ�:FA�r���W�L�y@�����3T�S�j�fL�?��w�R�m�<�@�s�S�Q�CR���b�|i2�_=��}�����c��}p|	����7I����Y�h}M���\rY�UL�n?_��`s%���5�uG�Er�5��Y�Ů;e�$^�	����,S����})��-�v�,s�I=��r�ww�A=��S��<�㉚:4p����{��۔���C��8���. �P���K�%����_���n$��{�2D��՞����^C&�ٰF�ܸK0d�+�������־�kbj�1���,X�I�=|�3m�e��`�~ຟZ$��[Gи �pW[`��,��Cdu7�(:P�a�@�`�����J��&ހ4)0(�w�M�m©%kL@��X���q�D��.��.Wb�m���T.�i�M���Q� ^�HJ�5 ������������4l	8��$��&����Q�$����\\�X��� *�Y��^�=[�p�:�mL&��N��
�
{��q6`Nq�g��S��1u [F`���L� T�E���u0C�w��z�N{d�i�F�d�ζ1��״p֐����	�e�|�)�怙�}���z1@�-�a�:�O�JW��m�'�Sy��$�	 �a��J�`�@�lE����ӛxl�`���వ5t_���7S.�ӿ�����2�~�Zv$��_[;���H#O���5�
���F�Q��t�J��F1_���p�ƹw<���2�Y�Rptu�-��=r#��J�e�f$	R^��z8h�	�=(q�(�2W0�:t�|Z�������;�����[�p��h ��"�(��lU�2-�E)D� j�N/c�b��N�f����,�-ѹ�g�x����W����S]M�y�[�AS���)$����ZL~,�}+ځ+���Rϧ�sQ�&M6f��O�;��?xw`-�� ^�o�|������p��S �� ���O�ȧ6@�U5@�P����TS�"�:��u=�]�ÌRV���
sC��5� /�3Aڍ�CI5��剮��m,Y=��- %�Q���������~+�������J�>��U�S�W.��#2���dV-ߡ<�� �1H�Y:�����Z�s% �.��Y���	���S��ӫ�j�
F]#r��B���'�F#��.z�@�B�<�l��=��tg?:��X�����J ,]Ȧ?�g�wб��Ȣ��`�6Q��	���l�f��=C�}+�����s��b�(\�P�X�V2&KF���!�� ��P$< � e֖`e; �(5q���UT���8e*��2�$�hG�Do�@/�hd@�a�	�U% Pt�]�y�L��&1��b��i<��z,+u����ıxp`��N�f�i_��zK�R�F���!��ȼ\2C9L�M�(-�A���:33_�%�J�Ϡ�l3OF6>�2�9���W�EVϨ���_6Fv��%�|��M��O������g	� nzh#<F�r8w�y�T�@����`�8�q,�
p���n�g���d�	|)�,��o9}t����=��P���1A�ʎ�m��p�2A^�t� .[*���ã�-�o�fc�1�� �j4�)�y���K����ӐR�]b�Vv,8}�T��,��M�7���]�wd�$[ݝ�� �;���q�<��i�EW�jX�4�d��۠%��!q�@SfL�����7	^);\��tV�'��[� ��h��M�4GP:��H.�@�^Pm8J��m�SAh7�)���]�a0:iـ"G
�_`��{�P��k��;��J3�5
|	=�TM����{���B�_�D����1�E� ���1j�X{�� ��u���0=++�V��Z�G�!D$$�.�lF�j}����'�������-z6�"r""<��TE@MA��Х*Ujh!X	D�H� %ҥ��J��tz	!����y��w���~a>��k��������.�����=u:>�����P9�/{�/�������H�'(�fd����~�U�W9Nf& e̜�Eq?\��A�4Z��AY��NpyW�7@�Y�(�V�^ѻ�hۭ����W�d�W��*y��Ӌ�vBw�~��?�o4�]p\��~��k=m���;m��E�oB7 �5�;��a�P�iM�����Rƙ�}Y�}��p?>��?f�����}���GO�(a��ҏ�tL!w�3��k�C���s��%��.��~��W,�z�l]�6p]�"3�ޓ�MR��s�g��w�4^����.�O5��y24]�ew�򛣯b�����5"��˳�'�F���ye3OV��m|3;*Rv� GEcPo���f�o�YK�_d�
6T�=�L�n,��#5]ܱZ'���5s�e�]t#��o<�����(�X=�u��^)~Q,'m֖ܞ+�����Կ��"�����9��_
f�/���W��uco!�?}�ނk��5��q�g7ll��@a����~�X��W"~�e�:����])���'.w`�bl��e�CfKF�w��Ա�,��&iXI�n��V�ցƳ����-����8�g���k�Ѵ��֝e��?±ԽlZy[H�rł�Ty��ԏ����-�icWA疙����6�M�A5�-����8ʵ6�N	��T���Q^�!�*������	��5�:��%ո�o��m��#���>�Fپ?7��,��Zߵ���D2S�p�+Ip�`�S<���W��wl%u�y�{.��.բ����UTs�(�ӏ�6�>�����y�3�Я��4|�X澝W�jpƓ�!VVY�'��/Dv����^c��3�	���h���cđ�������#=���.<� �ϾPf�m�P�s��|����%s[�T�G�T�;*0w�*��}�E�ܤ�7J��O����M1ph=�%���2ܵ��Zͦ�����$<'�^6�
(�h\�uֳ{�Ύ���u�f��k][9�}$�P,4
6y�~���~���	?��=�i�C��彺�����gV?��B����`ۉ2�Klg�E�ۙ�I��!˵��.z���=�d�n/*��Zq26���yn:/'�)���/�h����s+�c�~�J�}�t����@ɦ�x)��^z`g��x��>���myp)'���-�\Ph�����n�iY���v�7I�z�z�Aή����9�v�B,W�u��Sf�e��)������֓;��M	��vl%C��ȶ(���9x�o&($���$G��Qs�H	�x!t:;>���']��no�Ԣ�g����q��H돿�`�g�[���5���	����#/�ΐt0�V��h��LSu�^U��ɧ��Y�&�o&��-n�������^���ow&�^y:�j:���g� �|�{�`��|%
[?τ�?���J��}t79��^��o��@��)��צ���R3ٰ�>o������v���5�5��V�M�g�E�(^�`?�fs�d��BM�>����J�����N&��?'�%4�Z�&߽���&��,�{�/�;u�(���"y���o���L�X(#9��M<���(�@�.�2\o�;��V��3�}��wo�qa�׎ɧC��;�
Se����"��n�!)��uX�nAخ��N��Ɲ�e�/���"���)�t$�nab�iߥ�u-���:�~��Wϕ�EY� n\p����6��CI�j��[EZ��W��m�:eL	���������[�T@P����#M
+g���pG"�C�n�����r��$-lK��Is��n��S�	����|h�*�� ֞��e-	�9u=[�қ��ָ�e��Ql���	��7E'@�A�}���Irg��O4%�m�Z#�0�0�~s�'�@������I�f�F'�_;L���������A�W]0Y��g2�Q��z�f�Wpt}��˾��~��8?��3ek�:�M1�mk��^���ēj�H�����DfS�a~����Ej��z�!��ֿh����3۾�O[�����\�$��I�w�ϰ\�]ȡM�:)���4�]��RO4a,B��tS�NB�l��.٬����u��JY��G5�99@6IG�������F`v'h�,�/��b30*��2�������q��  uC���k6/�'��.�nD��=>��{V0hǄ�O���o�M�=+J�b�s��!��.�x:�M/�ϾO %�..9h��9-m�s�,R��H�e�����Ue҂2V�4,\X	��ȆC<�	{)�&-��j�j�1� X��D�ӄEV�	&��|�q��?�[�˖���v�CJ	����.�7��e{�)y����W�k4/E���� ���1�Ra�n�1`[7�uH���B�����?
�X�y��'ekz��Db��8��Y�j%�h4�Lj�e�G�A�3�Í�Ċo|Q��%g��QŇ�]���v��|�9�~�.�+�	񞼭o���EVőV�����fOCNp��CA6�BOhը_A�K���]ޛb�����l�5Ͷͥj��8P�?�/V�(�`7��+f���bjU��3j��*:��x��3�!�Ch�_�]���tuS��Y�B�"F?>X��@���w����d[,U�6�Ű5rowT�{3�416������
$��?"�/��M]�SMU ��7��W�Z_��:�6�$ح͙�P�2�.�`5F�kc�"D�f�g3qK/Q'��K���8�i���OYL�޿���5�'���]3R�ʱ��"���u�<�~O�ˡf� �L}��&g6�E��'��ܯ��g�� b�'��!�~w�W�V�N�����
K?���������S��S��z��J�[&��-������\��p\���K���A#eф�6�� ���/[M>u{h󾻒��A
�q����d�&����7�zsvc�f������̇�|ďWB!��L�E���F���LZ9��������|��3�����ցF�!�X���Ev���(kz�?�p�C7-U���跈�?哊�i��.��G��$'�s|2ȩ-cb��+��I�؉@i������)#E�{tӜ��꡵`���sJ)W��j8)p��z��BKJ�A���.)?Q@^ƿG�lw�ԏ����$�D��A���P'������9��D7`�^���R��J{y[��]W9�-=jͱ�6��L3ģ��Xt�-�)1�买�rP���.ю��/���4�6���gT?KB��38��=�����f�����^�ʪ�#�u�' R�ە�,o�@���{���o*B;�}W.���~g�ν �Y0~�-f���o�nI��x��7=i��-���;A�(0���b0���6����!��7y�5��bY�3���;~T���F�q)���HI����ߪ鱃��� M�QRF��rl�硧�[���&T {��Gy�+g��*�M��4�$`4J#��t����)2G��@uT=����=Fb�(
���6�rȍ���О����*d�F�����T]>�`�ހ�߷��\d1@�H̺"��wv����q�$/95�����ҥzC��'އ�"����]U�,�6���mllx�����-5}�D"p�^��#�fC!z�����ۛTY5B�|�Uy�J�rx�ǻ�h�*���^�]oy� �8��Owz>f�1��H�+��Rv���f5"��PP��O�$k,�7���J4�#���t�0�"O�� no̶Ԡ�4S�7V��7�?��hOnz�t	/�Y.�ڼ�%��eG��:��R��[hG��̝g	�����/IS??��uj&�q����ݨ�al)5a]P<y�X*�3��P��ؐ[�,��EK��<�g�ע8�n,Ǖ}��׆�T} {������V��������s���|{j�C�+��Y8�yK�s�tdb�JSC�q�5��IT�Pa�+�2S�$���q�A��oU.�ox(��܍^����i��m֥��<���e�7��{�_n��5[�)������W~��
X�����H� �y��k������95���Ȭ[$�-~/ͻ�����),7;.��y�Ӻc�f+Ո�"�ګ��[����-n��4�!6a�Z��%���-�Zķg��I�UZ���
�#�'�`�4���m�{�F�ꁦΕ���v�f�������6놭䟁r��/�����n]����@;�pd*���Y��p�xcEP�ܗB§����r��IIė߼�C�Pn�PSmcP��Z�����H���E�9V�i���X�P�����5n���w�OZ�wQ��7\��h�?��T�e��{�����Y���l�&���D���xOT�s��#=��(�E��QeKֲ�7�e�z��k�� -l�Z�)����d�G���F����l�Gm~8��*o�i	�D���E������'�k�tA��m��+�mJ��V�-qtj�����*W�}�֦�wMz��V����#I�$�֟b��(߯��c���jڃ��Ô0��:������� �՝��𥧿�yj˄�id��p��4o,ՠD�$w*��e�ZÅ�[R�^6=����� ���1i�
у��Of�e挾d]��j�0	���}L?����u5s�����4�(p�\8���=sbw�J5CG���i�5�?�yE�@h����VGQ��[�x�(�Mw zZc-�H+�P�A2}�>n���͞���w�_�׽I�4D{ܬ�'�#�[��h>��E @�,�?E��h�6S~�KLW��~��-� ���+�>�X���&�+K�23*_8�^�|̚^ďy�O�40�Ԧ�WL�4]x\�S�+�o�O BG��֯�EWV�%�r�Vs_8p�s�
�2D�/Ab�cI�Vo������|��&'���l����oL���D6/.�8 A�L�	�dQ�g����������j��U�5��+�y��}����m��[��^}P�I��j�4V�k�O�˜?���H��r�J�t�4
��dL�7� � ��1�qX�I�Eb�4ba��`�RBp����*u�6�9��܅E�����M9���O���7�&�9L>ɮi��D�� m�_��j�;=�D�Y`�S�n�7�*�D9ʪq��UD6<Hx�/E$3��~�T� �I�� ��A:?�m�KM"k01rDϝ���N2C��櫵���V�P����	p&�~:c���o�w��^�z�.�ɠC��#��CC�&us���	e~}ZܢM�~���"����� �c$'��G�a��v.�&5���W:Ow3q�Ȧ��_��9��|ɖ���EmAҴU������9p�� a �6��t�gi�v��YkA�/� ���]��˂mD�����ѩ�K�1���B��ؐ���Cw��e����QČ�G&��L�v�o#L�����1l&�=>�e�²|���0��X�)-݉9��2O	g�g���`k�4:9�/���o?Z��.�ى�?W�̎c���m�W_�뾁8T����m3����p��ߪP�H=�L2Ra,-'�߾E�N������[T�x���6Ќ��	�m4� ��w6�
fx#n*Y�
F��?���Eao�;H�d�ƌW*��ƨ17��K_B~MكKb���%7���oM���?3��NP��U  Q�*`�mY�tbPpG�����Fvȑ�tҊ���J��8~�;I˖mِc��t	�Z[�C��ǨT��5ʞl���g ���Ƈ��o4��?_���΁:������K8�(ٟ��,�ְ C��M��Ma�a$)�Mq�c��C5�4�`�SD�0��$o�XR��LE�!-K�0���� ��8-}S���D`�<7�{�_|^�07Pd���C}70$AY�Ugn�Ӫv>K7��}+򷲁�"ן��4�Y��`ZY�vM��t�("��rm�ʪ{��rL���y��&� �5%o @R�ay� #�PS���mJ���P╣�Y��G�ݨ�?d��YǷ`p�:
��J��M% ��S�m����e�w�~��LX�^��̂���dtwoT�	�������Юj� �b��Y��"t�0]��9���W�1�O�ۊ����JlE���E̓j��n�:���CFf���s�l����N�`w���]��[o�e�)�<h���I��q�W)ᮢٰ��cUm��}��k�R� ��d9�]0�0�ψ�u#d��R��9�R3�ʬ�kVI����^�N��UHD;� ����hY�8p�U^�W�*��W����H����13�͍=3��t��F5���$(UıΨ|/�X&���x#tf+\{�ՠ�`�Y{F�l`o�!Ur�����M�Z���s��*�-I!ݠ��QH��7�U^M�6VzH2h��%��z4M�k'�qc{ ��MX{�W�y����*����J�Y�.&�׫g~��B-ا;*���8&-2���ƈ��u���d����u"���h֖�k1�D�5�G�^��Z|�7�#�x�NBm"�i�����Z~�|�-b�Gy?l�kV���d�)��հζ�Y�����O��$'�sE�eam�#|�κRLB�^�o+����8	����発|�R��[?�U�ڒfۙpTmVۙ�2ȱY��e�}jm�$���oj��s���$�(�\tIm��f�V=O��x{��@6.�1kvw�m7a= ��Aݏz~B5�9:��4�R���;L����H	�'3��Z�3��@`��nw�]%6��(����v�(�q���`,hg����aj���+W�����/��1R��;:W� �̶��
eJ�$�Ąt����m�X'��~�<,ʂ�}�yS@:L#^�[9q���kk>��g� ���)b͹#:�g�%m��Z���׻�B��|94Z��3>��5(��]��&ɣ����}��&�HӉ`/�߷7J���k��Zqi�	�� &�޵}��eU����nE4������:�a���pE�	� �d�6.��2z��A�v�R�Vy P?��"	����A�|��&�LM���2��0�U�O�\P,�X�| [;��-l{�������'`��s4�}7+�\ɋ@�\�ơ�)�h��x*(�Q�h�2X(���#�D�����t�'L��&��r})�b�Ru7\����so�F�<Xm�s�c՞�f�s��T2�Ǯ�@�dm{�<?(����0��:�H���	����@;t#@{�s3�C
W�:ՅH?0��$򈱕~z���p�h�0X|��u�a��;}���h	T�8�~�]a~���!!���,�xQ�yWS��Z�j��Q���,� ]�z�aro1B�yP��E�ao�?ӡ�����^�;����4�(�5^>0` �U�)�q�?|�r��oajX-��QR~T#X�NK!n�ƒ<�P�'K�є�0~7 �Տ�مEN�QH!�\��O[+�_~��.���
r]i�O]=q�D`��!�M>�s*�Z���l������&߳O�?پ|S/�	���ĺu�Z�e!j��(�u�f�7�Ȣ������D��)��o��F�o�+H��Q$;Ԟ�i.�Jt�nq�� �F��x�!��֔W� D������QU��?6گд#�5g�Awo(�.�X(��t 3�-s���ɥH�_=��)�ƞ��wk�շ��j~Am�2�~�9��}�s�'u��ʴ&���6��L�j�qД ��'�����P�4F���k���RN���D`�s��~�Քq[�UeJ:u喗��Qa��]�:���&?����t��N����ɒ� �<�:��!��p�Wғ�S�y�wv�0b~��^��tf�u��ztƐR��>�Y�Y�fy��4�_x�l3F�`@hӸ��wu0��>�����y�N�+�����o[�W�pvب�@�U������ȳ�e>=�%�
�Rw[7�N�4�>t�R#�e�,��E���,y<u�{��V���(�JR�<VdsM0?*���b'X`*C�����r�R�ό����Ӱ��1y�PaN���԰�'YY5U���}���1�iG�);b�wf�1#8Y�Eͥ ڙ~���C�x�n��{�J`냘 ��8��Gb�xErۉ����u����M�� sn	N4�:n���͹�Z�ʃY��EW�Vyz��f�_ 8�R&K^��\~� �LC
�x%��7�{����ɚdk;�Ք~	��Q�SE&֩A����>;��Cx�L�#�?��43 ��9?�& �_����gbŌ����>�Za0i43��䮂R?R[�]�r��[Ul-"Mc�V'!�S#"f�X��W���r_{��D��Oޓ�:W["�)����5趲/�-.f�a�U�y�5xrD��@A�#Y���?y"J�#����\P�Poɪ�7�>@Ǖ�M��Zbn<7�5������
3�����qH~�ƭ�k%fw��u�8�~�E�/�.�� Tď�),X�*�ݑ�۵�(��w�o�pW{FƱ��� e�ƞ���M��(�x�+7��I�
�Xۜ=a�S�w�w��$0arR<T�nC6O;�"5��C馛�*����F�}�Խ�bZԣ�Cյ�)Yl��k`/���dq�7��>0���> h�#����M��F҃..�p�����=�XU�����d������ lo~��6I Z�1�2Ӟ�=}|uv[o��j�y:���HM�U<).��Z�s&��	::�x�~`�>��|���00`oW�+j��P�����N���kePM�`���u�{�a�_U��4��mϏy ��Dhd�fط�s&��`wҲ���_�ح� .  @ ��Z���9�SY�麄H5�\\�u�gf���V�E��ؕ�ULn�3ۤ��1�V@�U�K��m�L~����@�p1:�Z��J�=�'-X&C�+L1�K�������a�z�~5
�����E�4�)��T�Ct����geVʋ�j�J�>HO-Ϟ��n��ܬ��x\�J�����H$U�̓�����>�r����[xjmQ�� 8@�*�h�
(m@g���jһ�+Y �e�OjGdrb��,c�]���M�[m@�]-�����#����(*=�,= (��XFJ(�Y�Q�9��}>7�	0�s.���؜���I�;�!˓���G�k��C��E�ڛ�O#�w���D*#xJ��1S�K�)OM�9͝�~[�z�cfߞ��k�qvP�����0��̨�T>��zd|� ���T�wv<,�b�=<�U�ph�u&���i(2�h�%�D�2K��7�����!�WXF�l9'a�r�͑vy��rL���bc���|b�	�q2C X�
���`�ʦu��T����i{�������$n&���sc��̀>��X�hS�8��(�L�[��W���H�g~�KB(������˻�Ӽ��6�E�~	l��&"�H�{�B�1�LݼzRWM��əFȲ[6�Z���fW����+@QE���"'��D1��c#\h{C0���?����'��@����EU�P�A�ĭ�'7����mx�dFGR#��6�+�}�-��1�ǘH=><��A�T׭(���cyӉ.0�ת�a�&>�,�����ۛxt�5f��Td�p��=(�rS��c�T�J&���[�HM��$��s���?WpLҫo��D��)�fˍ	!����l���^v��MTg��!c%�a�AJ�jO� 	��o�R�԰��ⵙO?�(~�/!3`Y}�� 'S.�*F�&yZ{_Y.��G�J���Y���=oY���2����'��{~Z�yS�{`V#��-�Y��"sn�&��G�S��6 ���<3N͆�v @��k��obůtЧ5��!�v���#;4� ���ß ϕk��q����d����s�;���M��A��<(�h�[85k|���1�}����*��k�)��jF��m/1����FYA�K%�����So&f f'�a���gҹ&�V[�4����Y�SI ���������C�l��xo��jb�^��V�+��y����2FN`JV��^O#�#��Y�!b� t�o`�����>k&|���1x�א;`y����b�$o��]fc��<�s���Yj$�4|ߕ��r�/.pTO]�M�/�a13}�M�a}�k�0ݏ+�{Z��[�Ӆ��CK��Ͳ&��"�N ����d&Mւj�Ԓ)<��͂��ՇK��_�QTZ�4���^i�aL,��|W���,������ H-��b� ���c��KwʏsJ��e����*��~�1���i=(V�}/fϏxE!\�����r�{�"�+/��N�%4H��x���Е�V������F*&x��m��b_Uw�OGv�ږC��VV2ˑ�>m;�(|#9\��A��kJ*��j�0UA�$�h�?�
�1풐f����#͸�g�)k���<�?��D�q�ӞC�#Uբ�1���*����=Wf�*g�[R i�9��S���%��� �[����WI�����z�3����Q���7;�K՛�u�<;�����̂G���ɚ���e�_K�K�Ʒɥ��|	=|fu[��%*q�P6��n��l |���U�Q��2ﲇL��I�lwF@�M(��5~vVm��]S��S����_g} Rg�j�;+C܃F�V��qo�w�e�F��L��B�|uN���g7#H	��  aT,,dw��p�|�PB�M�M�9��pIh7��I�F���/ ��w 8�ʊ�f�H|x2P��*%*2j:r!�4��d�4�$��Yj%��.�~)�&CI���7����k)%���5������~�w��^�����8�W�90�R�]��3s�9��=��fl²��w�cfR���F��s��k�j}R||c/���U6(�2O<H���}��n~�CYI=��h��Z8J_�Kj�'Ƨ^<�$�����0�Ң���)�8�K��[>{��<�ln,���yR��K��Cϒka<�P��d�u�<R�D��O���[��h]Y~�u?]8]��	������f����QR��⚨��a~ڇ��w��Z��brI��S�\"�n1B�����
��ky �~X0vƬ:����ڻr��L�x�+(ͻ���
���״����ghl�Ҷ����=�,=�+&�Q��,�r{�D1�iLoi�lʐ�(qݮZ��T�1�����ni&�{Y�#���2ն���| ���K���݆^Aȥ3�3��
�su"~zN�ZLE��{�E.��f���X��K�;��=�/2po���v=����s����CЋ�;��ܽ,�*����~恮�,�-/��s���k_U:O&O����/�|�sa���v��G��Y-��7��0?B���a�C�:vH>�(u��[�����ۥ����u���j��߰��bP&��s�<���oWI�T�<$�����h�8�Rּ�畻�b�����L�t�:��_�$�T��3̟/m޿�@����&��!�[Ԥ�I���_Ȕf������۔�Es�ci\���j���J�zS�����O˲ ��'8��Q1ٓr����� �^�]|^9�ss(���n}Z��*��r_RCd[�.ޣ�̳W"�J��_3;;%��:��fI���鰍��@9�D"F
o
�e���|8k]��].����)PtKI�A�C�9p���d.��ioN�I�����Ç2����6��o�VQF(�]��zU[}�}��m쉣Y������s���S���j���YD#oT�Jg��l���*���4��%5U1����)� �˾x"�b�DGߕ�.#���n2@J���â6�f��Deg;!�������x����WE��/p�{��)q*O�o�Z�}h�P��4����O��Lƛ����	N�u�Mk]���G�ĩ��m���X��@n�Xմuv}/�A��� A�}E�lg�:��h�Y�_g���2�9���lWP,�"����v
���=
����Kg�������j��]M��	H���a����mCu��4\f�<%v�f�9ծj��>�#E�Tw��?-褤��_�������������yc��J�7�;��Vx��J�f~JhH���_��6�s.vӁw���4�I���y7JMw�R��u  QVg�.������`�G�U�n�����e���c;���_�n0ߟ�Ϭл1'qR'e�dTW���nT������K��kx��oU��qB�x�KY�2�E������N�,S̵ت�C蔏'A1�NƛS�:��a�\;V �5��±�YFl*�����{����2�/�DmhP
���I�,�y�ª�*�`o>-��~�#l�t�Hd��RX_ݕ�K��U���3�2�ʌv-6D��||:R��͋68'}eK�P�+z>�uCB�G"��-��:��Œ�!R�boK@6k�� �ݾ3�~W>��e��Y����2�#��a���`p��'�$k�dɷ�v�-d��k������|��l߿���o�'�ϱ���Y<�S�K�^���׉s���S�W��ߔ���X�@����}>��DX�
�u�TS'�m��6����B���f��[�ٮ1_��=����7,�<�zi�}aM��b�=�k�[~���}�� �:�>y/�������*h�,��!9heh�{J����7Ko~���Q��/9,�F�#��>��i�dz��vc�٤�⥃k\��ϏL�ǖ��1ȘYK}fR��5�����G�}⭆��J�	J�0��*F�}�����n0���Ȥ��KM콢mKC�C�T��J��ڬ���|W̫�m����δ{|Ot89� ��Z\H����)Y|,���l��d@�͝M�(jŒ9��i�'��.{_og$�ta���c�׬���݈��Abe���g�W'�����S�Z���	��"���-s?u�"�e�f��s�ՈOj7�i��NTF��-UL����ї�.��s����;E5nl1w� �F���[��a�����RK/m3'���f��� �)�UtUw���=�C�9j?�Fy�\{�_��N=�$`�@��h������>OВ�E���+Ay��a���&�2o
	�p�	��I����R��?��������.����g9[��]�v�d�[��n��A�#E\����|�}~50gQ�xnq!�P�B��䘿��sP��p%�dGM���h��y�9�3��j+ȶKJ1�Ė*��J��Mp@��p)x�I��Ĩ��s�b��\Z"�fӛ!�cja�ףЊ���ǘ��jwY�Bu���
3�+>r�������8m��B�z^Lg�Y�wߙ��vE7a�E�'p/��<~=d�
+�Z
�
��}<8��ԉE��#\�h{aD>�$usz�ٷ�v7�����_�U�ӷח�^����K
��+���.`;}�*�pB�U�BPø����m�
�S[��3�P\��H�?�n��3�T��z���Z�^��o�p�n�/�ϓ��I��^Ξ䎾�|~�����&���XEX���Wu8��)���wR��W=������330ҫ�R�Ng67����m<�y-z~�`�H���dS��,J�t�su�V>x��h���jn�x�rA�����C﷥���zw�W,�"|ld��_�6��]�2��fg�2g���0\&�zU�*�SY>�&;���q��T�S��3�w]U ��iͻ��.��c;,�����ZT$lpKT�_����_��8[�Z�wd7.�<=����D���dޅ���B�?`|%�%�F��P̑�<6�յ�~BJ�b,���D
��";:=���K�#p��DjQ]��g�_��v�	�C�j�>#�g��u��澋�$W��x�vZ��Nԓ���c������t�� �`Q����ߺ
��^dW?��S1��;�=�@��_�g����i��%6'�p�ؿ�R����S�-�� �~^�q�r�f�d�Ns�9qG�У���Dx���Z�����PK   tb�X��"�IY eY /   images/8cf56d13-717b-4162-83ff-adbc9fee247e.png��e\�-��{p[ ��[ �\	������%��,w����^������ef��7�5]]uΩ�0%i4d"d  �&+#� @�  �lD���������@��!  �J��0<1@� јUw���� �~��A�,炳�W9���O䧂;>���o�~������*�j5#O��y��Zm���|)�i��;��׷�9>�^r����y?������|�
\=����d��ִ�ԇ��Ȍ�l Ix~���6�(``i��@��e�4b�-��\�N��wBS����"D�^���_ku�a�H�c��ΟK�_�wYC�Ѻp���8��& I���5�aǵ{�޴���b��l�/����䍚Ԋ��ޒ�aÖ�¨�w��Ce�R���r�AüE�Wq�������D�L�����mImkI���w����c�}m��à��r��?�;�{~��IRB�'uϔ��4�7��M��+G箷d^&Y;����_&C�'�Vk�4�f��o[q�(E�����5j#��a���ލoI�����jȓJ�	W���k���$F��v�մ���5R魍�˝�\�M�N��VK��+�>��18���Uw�۵�d�f�O�_���<.��k˭G��9�[���w�U�4�ԲM�py��A}�U
?xP��rP�(;p�-J#��銖 �ixLD#=A3~�|C4���j�*!Ǆ#��y���7��v�K�#��G��\���� �4���B�8�A,����R��@�	�<Sj���qW�|���)6��
G�fW�&gL���-/��-M�D4���"�(��@�u�hD#B,�2��F~�-Mo��×}j���n�e��F�
9�y��rPL�"@�*4vO����1�̲)��;9v<��s%�M�|�.�.f�*b��j3���al͋�58�Խh���L.���*�����Q9�S������-�l�t���D��6���.�A,6�����z�_X >j!B��!�Vxܛ�&A��V�ˋ�*V��~U��G��1q��9l�Q�"6.��Xg��_��;�6Ԛ|Jȉ��m�ұ��;�N^?<n�>��&sb���-�����������Iչ?S�=]�V�y�w6�ԍ��(e�d���`��6^%Wo(�]���k�V�E�����E����ңm?��-û#\ٸ �>�}�����q�����/}WxA>ҏQ�~���$9v7��4����D�h{{P�%v�ۿ������o�-k�_�8����<f�h����̶�(}܁ ��$-��#�S/�.w\�way��O�^��Bl���[O=N]��c��?��H�`GͿ�����d�b_m����J3�V�_����1O�%���O��:]>kj����)��	6� 9��h�~�,�~���Խ�q��|m�̙='�T?�-"����dV�-��M�G��,�'�8׊<
-����^�%�	<�V����J��׿�gO������������/r��[U����8�$�cLf{�兒���_$]G@�H:�Gm5\ݜ���
�&*9Ǿݟ��r6�rKu�TNڤ�>�%����jA�\:�������R��Ф�|F��ᝥtx�G0fAo 8�M�����僰_�F��s_�b�Q.�'X-��
������/����E&�,�;��ʀ|����S�ѹٗm��&�I��d�kE{ι%�����*S�|��: �a��O@I�s�s��Sҵv�j��b����O縉�s�\�z���C[�%׊���kL�����������|�%����B��O���d���˰d4�:���⢎R�e�������.�[A"���e��?
��
L��Z�?�{8�����l��%��R<e-�Bu�0���z`~�]b^�E�����vhE��{9�m��y�nϩ%�-���N��y�}C���&�T��ӍBw�*��ȇ�`2�6&H�+Z� y�á����y�"^��e_z����s*k͖��U�5����G'4�NP���L�;�����<֯o������q��W�"Գ�l`O`�G��q�b.����9b�K�zx�]��r��a�V��}Z�z�Զ�ZC_$����f6n�GZa:�9jQ�	�$[�GE}��[�������� f��MRӃ_c?��y`�C� ���/�3�2eg'�Z^���mob�xH��E�WD��3Y��y'�l$1�Z�h�m�4F3G��RQ���OO��u���Y��n/Pl��A�X_H�]�m�����>��?��/@����Z-3P�%�̯uRk�T�H�����P8y`���Ca�[�ZP^~TJ궴�Ǥ}aY��D<o�H���t�nr#1�Q���'�q FRۍ���QX}.>'�g��R��h�)�-^�739��'6_M��
����tjez��`ԡQc 
H)Ň`�k�<�� a��On�D�,������o�^܊8�㈃�#��b��a�k@cї����S������]ZQ�qYڬ�h�u��|�}�~�@[��}iފ,���V�q<�D9L�B�y��D`�#:j�͊�@0���m�ș�.��K�����z1���� z�m��n�b��\�� !_P���aM�)6�!X�pJ�.����{��3n���/ʲE�J�Y��W�_�L�d�h��,O����=��@E��2��h�2{��AקL��V��bf�Z�?��Y�����\�;;J�lw�\�<\ќ�L�+z���0 َ��)��$�S?�n`��lW��m��M���@�g�����f��o;J�6��������5X��뻈���t{�v�p�B��Ll��+7lkD�\O.E?�6��|�a5�dZK������]��@}���EI��/�9qk��N@o�Y$
es��I�+F�����U4K��-	��c�w���~�X�����cM��:��ή
v^>�j"��<�Y:�������l��5,cf-`b��ǭԯk����)ÎM�dZ�F*-{�X@ɹ�Vju�Gg��"˓DU��W�0����k���Y���.������Be�����?:T�O�VI���OOO��������U��.�W�q//
�uu��WTD�t�S�	�����|�eH�s-����/�4��ٽ�V�y����6��c����e�&qt]���xy�%yZN����S��`ՙRC�O�ޟ�ó�C�3���ܾ�Z�Vepۢ�q�"��<RYnUt�ν�v7��u�x.����m�Ε����W;�Ț\���%L�����몫I��z�"�ك�77��(F04p}��Z���}?�ՖX�d��mɉ�*�:�����*�:leאs	�up�5����R��/q��WZ�&��^�\SYUQ!S�h۩SRe=�ۣ�޿���Ȱg��Fۻ�~���l����T��.�5���̧M�v�msZc���7ww�G�Xb�J�r�G��IwK��l �Ӯ�3��('c��F�Q<��(^�ۣ��y��Fk�U�۔�jy�� �X�^��xb���h��"�|������b���9�s����n�fT~yu�U)��5�?(�\}�����RÞo�#m\T����c2�ƟN]ݱC�	��Y7������y������� �
S��RL0
TL!>��6�ɱ�0w�J@l3�in�u>U�4	�A"rwʗ�	�P���ԙ-d��T��/��$|��	��k_>0����_��'�u�'�ؐaZ
Y�ۧ{�3�f��O�M,�k�����8??��Uk����~�gd<z�,E�:�Z������~kV�����%�k�>[��F���¶09JS�@��&W��A����x�2��=z���8�*��8<�Z����7�C��J��%oE0$v!?N�܆���"DtxVw�t��V\�~�z�׿u�����+6|��=Zq��P^\K����>30Q
��F��ۭ��7�I���da-:VG��e-�˒�kv��,��B���}	<�'m�`������)�땏�y^}�:�i�>��?���Z���w�'��#�T7��tT.'�m�O�i������~�Ͽ���ۧ�~ ��2���b �E4��?ؤ���[$�>��#|�d C�w��P K�$��*�s��7�	�._�®��:�0Q�8ax����D�j�*T������!�Ժ��������6�]EE{W���mH��Q 8��F;!�V
�dv�?U��T(�����z���:��3B�d�G5�==I���7j��zK����/�p[��uJj�z��^��d��XdRe�m���J@��a$�7b.�ϑ�!��%/W`Nd��B~]Vշȹp `�����~�`"���)�_O���MF肠�,k�h�a��x`������N�"�+�bΩ
pQ�KR<բ�<��o/��SF���J�X��4-ɍ[�{��A�]?V�0���H����i�4��|����)pY��Q�"703~��\>�/�\NI`d=oa�-OO�F8��t��D�9�<�'S��܆��8y��=�=f�#hy�|M�뮁��k���R�VL7���`lM���}2��!=�n�?��ΜH�繁���2uf�o����$��/eJ�n�!z,v�G0nok� $�ew�c�5#���ikˉ���Ŵ-3I�ihR�h릢Q���%�3`"�B�DD[������a�|T�%r������+W��Wօc@�����8z�N�G��G�**ܡ��.�'��-ϛ�(���d���
�Oo�0�����k��+��8*��e4��nZ	r��a-�T��������{?��z�o�a!��sB`+�|�Z�pů��r�1(*�2n���N�}�W������_�R�q,V���,�R���ItzȠ���]��0Y�*S���hBw�/��|�*sn����y�C����B:�Ym.Ϣ��o�!
MLA鉨�CՆ�L�� X��pۚ �F`�w��06������_�Z:FI�Y謨v�_Y�c��n1��ϡб}b�GĴQ[��~����^���)S����|��/:������q]:� 7*eFD���������<�r
�����v��u[=]hu>X�]i��[���R�q�z�C�����l�����J�<v9��h���@��q��r:���'0mN��ʯq���أL�K��Y)09&G��wd��8�Uw늳0��!bC����)BT+|��u);[�j��1`� ��&tNW�I��62΀��@WEV܈'�d:�b�xּS�$`y�������B�QBj���J�Ť�T�Ч>A}��Ak��>����7,,h£CIg��	���³_��R�06���"�WO�"Ʉ' �$A}��	���\�p��[o	deeƫ�<	W`���##FDM����C���ȏ������wS��s}��Y���z�7��i6g&AYd�	l;�����S)���_��2Ca@��O�Y?���ɸ��ƫ��r��+�)�|��m�~��JG���Ƴ#8�c�{F��h�rܯ��c8�#�k挒�t��$0b\�@�v�����8
.݃�Xwā$��ǋϵ�3�.�L�3�|���]\h���C�(9@�N��n��q��X=d��&�;:��F�V1��u��,��rB�/1�t߾wm����U�(�}��$-坴�jw�pk�Q�J��jl�o��Viяk��$Fxm�M�]�H������r�}Y��oP�G���
��iEjof��'U���[����6¤
ڻ/ (.���W�0X��x����4�	$�IH0��o:Deკ�t��u��%�o+�ԣf��d�(���X+�ˤ��~�<�n�q$?���|��(��^s����Ӳ^�}��o�=��^5v>A�t���F� ���EC� R	���+SZ�"��+�_H�%͢g�@Y�����G�:5�g9�:���k@k��G�:K��.檡��'p���(�pj38辕��J��o�+������������>8�: ���n��=��<�O]�L��}��i0��`~��7���؞�/����چxp�?Zਔ:���� ih+��0I��R@��5K������yɪ]{�3<�f�:KN-s�U������5�r�P���'��ŸhK�i�x�ҹd�>���U�R�g�1�qۦ�i���s����P=�e���c�V�kO�읤FU�w�@�Cڂ�;���!��> ��P��'�"��I�@�<3�JyJ�Q0e!�3��$HD�$L�� ����Y�����(a1���;�Yn�&�A<��^?��]ݦ��,��L=�5�|9ЂOS�#L~АQ%��~-d������C��5F80�`���a끏��핎�W �R�v;��n�^EN�s���Z�����l"L9�9 �,��cWrw]�yk��i���27/��{�H�s�ְ��8_��
1�?+>�Xu����A{s\<��m�|RJShQ2����<ؾ4���
�7A�
���Q���A�YX�P5��Q8���/@Ze___Q&Ǿ��R�C^���RU}�]I�o~ïUC8�p[��"��Rə��N��;8І�郋�,��Sռ{�,��^_D-��$�FU��2�>�����UQ$x�]@�Դ��V��v��bU��#O2�o�����?�j���Q�.$C��l�u��c��7e�|�9�:ϯK���S���AY��
a ȧ�k�Q,c���^�_6��D�����D�f���UPqX`!��1��!jF��yd�T�>�������l1�xy~�~�ە��.�."!��A�ޮ�5�pG�ؒc�7&<��1v���#�4˳�����~_��!��������U@��yT���c��K��,�s� �|�0�{���ֺ���~B?[ȬiS��cҾ��{���� ���75#Ŕ�Ւ�h��HOq8ڴ�Y���5�5?A��xS+�5�1��<���9�O�gW����r]'E#x���c͡a֨����Y��E$�;L��e����eꙛ|��L�p�/���F�Ij��ڝY����d���(>ٖ�����(���3�?C��?cr�2p��H�m.v_���7�y.[w�����˺���gw4�u��������W�a�Tq~�`���y�%�0��	l��5d�����Ǆv�/�f+,�>vf�i�BW�!�Φ��V����@pK����a����P���(�h�c��,��A�L�)�mε��<nKU��>��訍�(�3�=Dp��Z�F����z>K��0�Ц��L ��Q���-WCug�B�y ��rt��j�bmqh�#��U�h�*�oo7�������mΣ�G��qJ�u:�N��v�L2��	6{���il���:�t�?�c&LS�
#(���9�׮:R+�j� "푯��&s��2�O{#�}g
e�|�36^�ls��ը6&Xk��"[��Ğ�]@��C_(��M!#l���L:N:��I�զv+��9sSMwޮJ>�k@�"4nE����]���4�f�Z�&og~����;��!J�W�خ�|��[��@ ����+F�����nJ��`�<�a�rm�3 ��J�ޮ��>J
��)$y�a�ǩ�s����ؤѭ_�Y׼ţ��b����S�VMlU��ʲֳ#Y��|�$�d�n��bj>�VS��K� #�?����%N��+�����)V+$�R�5������]�������,�W{������G�"��u~�����5��*񐲡���=b��j;N�:�#$	��֋�G��!!�9�Z�Y n�`ic$�r�܉��p�D���(������G|�6�KJI��edI�^A�4�|�i2������jI6��;���c4z�3>Q��+s�/��Q>�a]����T��FT��+$���F����&m�1�U���ٯ^g����Tc0s.�۹[���X���}[̹�@=�/�^L�.�sW� q� ���6�2�P b�|�������`����{�j��2L����T1���c��ߞ"��n��}��,��Q�b����UC�A���z�H� ֊����me#��	����P�Χ��E���
��A��t6e\L��h��:h�Ԅ�P���N 	�$��#z(�m,X��ͤ��J����x>�
%���K1z�H����~`1����=�Kȼ?����?-r"��x���En���8'EG�Z�������{�K,�6����aƨ���3ڥ���6~�����T��rT1
s���l��6)��I�q,���*Ċ�WZ�$����~�T@�ڷTs���~�X�k+���`S4�kϚo #I;r�iV�~ޕa�����
FàG�c_\j��F�!�_�Wt�U�1��c�?����KZ��ᴦ�u�p�9�r�f}/��d�3�$����J%����e�+��?tE��V膇����x�a �@*ꈌ�R^C��ݖ���h�։u�����;��c
]5ARD@!��<����u��<Py�m�u�ά@,a�X9�7�������w�E�?��xf�\��1?��vX�P�V=�K�܍�kN���Ӄ0���L��.�1j"���lvJc˖�"�%X�>�~;3�f>��.�+��Q��5���u�h�ӷ���PL��g\F�L�e�Q#'}�界ru��X�jn�Tac=hw�o��g�Ii�
ì�L���ўK0�$@o�������X�#�K
����e���C�B�=�H�M�ύ~A���ym�b0o��*�i�(�K�1ӊ��������U�/~ͼ8�/�?ԓv��Rם�u���w!O��*ΝM��p��⭮�靔���?�Iq��N��\Mŧ������6�O��q�a������`�|��:��tVi@�+�HI �s�)�˘F�{2
$�lE��Q1�\\}�e[ۢsv�N�ug,��(�T��
�i�ޯ��Z8"���G�9�������m� ���-�g����llV>��U��E��x4����Aq37��D~P�پc��^��v�֦�\��u�`"�>�Ľ67�o	�j>��t�[0⃡�d����8'_F2���*o��B'��npX���eٝ���|b���l�7O����ҰY��3���e\����aԗ��<' �}�$>�9�Ͱ�����Ԍ��FDD.I���jo���B`�ˁ!|������^F/#`O��.f�LCwr��t�#�Ӄ���O���Yq�vK�crI��}���l�:���NEv6�,M�ǻ���*��fb}�0L����V�	^���yu�&���g�!����������$	��Ws��|�Q��|���p��[E�@X����?6�c��3����Z�������nO�/4w�$.�d��ג�p�9�⩛5�"�4apo�ఔ`�	4�cJm���?==�(��%R��ҾO���k� w$n{^�H��c�R}�Ȅy�9�5��j�UBs'/Čb�\-}��|���ً�*Ϛڱ�y
8�06��,;�EW���d�[�~�����.����b��^��b��{�;�X9���d;ޝ�V#�(���UxF�C�N�ǂH��ʵ�o����\���2+��ջj����|�닞¬Ь#�D6<��i����b�ϋ��e~fWsQ��K��\3KK�j��m�04�H�	���].U�v�m_��JK����b9#dPi��9CԴ�^_E��Q�ժ^���tdG�w�hp]��bs�lѦBU��)��>�C:��U�;Ξ�YWw���گC�phёO�ˋ�~�(+O"���誫�|�!�+�p��y�GyT��/����^u�l���l8��Q�˓������{�C��\$�M����`,3l���	��Ήv�엻m��P��KE��*�h�*���`�����(j��)(�kK��kMc�-�<�_�c����F�e�-�;�E��N��Hٷ�#K./����7�����!g� T豟��]�4���m.���%������֐}/���=��*Y~q�<�Xu���gE�Bu���(C���Y+!o��������sSz���+��a��ٲx;,�@3G�r��^{\u7��n�4��""X����V�pd3Ič�!r0p�+S�綘�<'w�7/RP�St#9(^XX�8�7��b��k��naZ���^�ZKa�
�hhEA����'����J��`pB;�B�\FY@�����翄c��s�۔ظ�p1����Y�&�o]\��h�6K_�S&ĸ����Þ�� �xqE��z���l>mҵ��q����P�������+++�J��7��ө�j�}-,n4~k��N�m�d[cC���3>U����Ku�]����L ���h�\���jݾ��i�E�+�6�7�dH�=���#tJϽ4�yL,X�N��|�K0a�1)F��ql���M#Q�YhsԨbkC�F����t�W�l~�UM뺡�f������F���ea�m�Ŕ(�F�g�]�7F[q`(5%b�]0Ůu�C���At}��Ԅ�BмM `$���O,��R�n��)<��F�^��1BWC���'���v�Ĳ/�W[��~k�ʬ9�Ԯp��3e)-%�Uh">�]�!���|e�J/w�`��%��*��p���g>�j;�!%M)̄uh#3ޡT��1VF}�ko�@��-���w��w�$�d�|�xS۾Z�QJ�B2�0P_�`�U����g�Np�����7b��7��y]#���/�4wޭ%�(�_O6�rs�Fr�o�ttN|�%�f�קb-#_��r�����%.��r��Mg�~�G8��)�ܒR��V1��{cҤ$�\G��ߛt��رg����f��%R��*J�[�fY�i�`�A3ԤN�f�
k���N7�ߣ�@�]&�-�^ɮ����^�ֲO(/��	���"�%��y�:�6����C�v+��k�wȴ�3��iM�������b��S�*���*<�j��b��V[\\��-������#[k�o�$%�@�����;�Y���ş��N�Yd��/��l��@�@��ގ0N�>3̻@m�ņ!����]�֐9C����B�P�7��C)�+��&��p�l=�\��:B��p��/�|���[_l]{6��L�B�C����W���?0�eWz�\t��8�/]�eC�t$Y�cz�����D���7sUo��|��:�2��@2��������wל@�1'ܯ$lK�����4�$`ocߌ�!6�di����"�E,C��s����^�@�;�m=�~b9��3�w�i�)m�#3�Nu@�����u@N��V�KcO{��+�<��#|�p��ܱm�%�~�Q��.9ܑE{=ɽvq��4��ց�#�P�X����vaF�u8�����J;�Mk{YDȕ�{��P�JC���L SX0�P��`�����G\4.���A��U)7(�9c~Vy5�h�4�+�'��M9ZWz��Ԍ���A_�����*�6�a�$Jj�� ߘv��.�����`]�Ѐ<k�J�������V@v8��X�c9���`M'���A=��ں`BKH�e/`�d�]0k�����S�hZr���`�����R%ȁg���B��Tl�$n�������K�@�rߍ�n�Y�����ɶ0�LA�I~pe^�Bw�I�ZG'�'�0H0��:�N5�u�Jh	�Ĩ��5�c3���M��lL��=�[�MY`�����q���gDu��p�A1��:S��2�|"z�4ݦ���ɘ/��,�Ҩ4�%t���S�$�LO�Q>B3�NL��2_;U����=7֞������&/���i9U�a�x������"8�Foc�caEޠ�i�
X�a�v�x�]����O�5g~1�i�+�zk����FD��r�qD����p3���i^��N����� �����&�S��[n�S5�H�5ĒJ;+�"� ��g�����B��荋x�?��J�bC׋P�+�o�#c]!n"\
Kɚ�T�
�6�i�3��p�\}�פ�a���O��Ltg�D���-ͨ��w�,���2�W���P~j��$�N�vsu�PpN▹�PO-l(G�Ƿ��r��mQf�a�=]C��_$4&1�� �Dܨ�(qqѸ~�)��:0���E$��ZK�����|LL�}&@ս<?����+���?��A�|
Ke�):�O�c7_ ƹ�x;��4�� �BĞ�t��?���]M]�����/ bs��O8�����5�P���J��GnifY!���j!&"zr�&�5�<=�Ԃ�
�ISx������pa&�G������
uGG��	Zv�����ȳ�*�^��RB�Z�.�j�D��f�n	F!1�֝�3e���@VK�Dێ�Bl �@��^h�ց	��fw�bJ�4.��晌p����ٷr4jm�{��('�'�7���@��G°��Z��q+ip����%����Lm^� 1��ZDQO$"/���(΂��j�.d%@�aW���8��Y��v.��Kc�����>.�g�ܐ=�ְ�����&��5\k�
��}^�szB�9�P�UK��t4�s�����c8xg���RX̰�3X~���o�\[��ԶT�v����y�t�y��;�5�1b(G(�mB��K�7x�c/�X����ʎUP�++%l�|�NҨH8َ/Aǫ��~��e��H�,�A�׽�i�#J1�C$2�,$+�Q�@������T':V����$R�tZ����yђ,���Ԟԟ���|�c������'���F�{�wk���7�#�5 ���Gb3����i�DbwG��v_��~FI��TlߜA#�`ґ	��A�IҎ�3���O(��]'!p���g� "U�`1\�P��eu�	m�F�~�ʨ�;Z��vDG��B�޳"�ˀ ����E��4�_��U1�o~��65���{u�E��]�8�HD~��<�����oGycm�2�?9�!B�k����%6�,,h���8�?L�ZB9��ؽ�z�I����|0�j~��ށ:�TjR2ѽwR ��(��bր6�X��TD^;�Q S�V�i�V���~��l	�C�@�>~��Ȁ�қ�uDo:M��V��+�SKL��a��l�hQ9狅<��x�)8��d3�XXrhY�G���%��[֢�G�F���"�t�ON��)�S�5sX��db컗�������|��ɔ�����59�ސ�b�HJ�4�*Ej<���r��:���:��Vr�)F~i��q\u�F+��s�_�/�rN��U���K2'��2��������.�N�"���;��U�
%��T��v,�}�i&)n[�o7%��2A����r���#�P#���}h��4�%���'��P)��)p��@�Ts#�^8�st^��Z�����)�CE_u�J��E?�+cDTJc�QO4
�-����w��,T�2�;��R<���;W��/o����"�e��Ʉ?=t� '�SH:�O1��pjK��L��P�ۣ	eCI2�2��w�$�6â�T�H�cB��O�j���X�>���S����f0���sh���7���	��;���(5���?���/���3�ny��_σ,��4��
���׻eN)��3�6����n��ARw�����H�I�w� V?�4qJGI���SZ�T���������m�O�J����W{���<�+�<�C�?t�Z�AIA�3� 6�����PRb��C��j�W3� կ"a[}�lLKl75�'?��Y��u7w���;�}m��fy_��i�P��3AwH��/��Fw����18��C/zyX�u� � ��c�@���¼�E��ge_)�5���>�@ �a�%?��<��!�8	ikcc�Ņ�_Z�V*���:c��@�އ�4�A�D��%-!U`G	Zw���Y�I����8Y���3���p���!�,�T��獛�>�z�R��0��D���FN�����l>GJ�_��?�n
�kY
�5��|O-)~���!�7}C��HD��0��q1>��I�+�!�Yl����,���LMƭ��8�Bq�Lxb�L����]ꐕφ���|q��'��S{�c�P�׿�����EEu���8v�z�Ν�9�����Lς�_����ȝ7W(nC�z�����.�� �8l`
����yw�4�2k�P�NQQq,��
�����#-G����� �[�3���\�Ԋ�/2����c��gp�>�V����]@�
A�#A	�����^g�Y�-���F�Ʒ���GrlyC�!6���U_��`���Mafm:3��*o�܁����v��q8�����yVV35�}}��Wڢ]���S�����P�x0
r����~�ҍٔ���+� `K=�x�[p���Bz]�x�@�d�V �! �M�	��X���n͈i���A���E6�-�a"pH���cGB���1���L (�@
DS�.��t�Bt��5u������h�ll@z��;�h�����d�Z�_Ƅ��0�t��?ȁIWQ0�l�a�J���.�*�%���Hl0q���
�����!�Uua��S\��сDJ�����	?�&
a��t��n�No�y�<"$) �&��~	�.�ͧ:�	�f,�]�旇�Ů;�豶���z˸O�*���EG���?m����Pb���ƣz��<�� w=�BҒڀj��c#u{H�
��K��(Ky�)�6{(ߖl6dO1K(���d6f�|�>��r�e� ���B�}��4&��ڃ�4X[o1�w��g�.�A-�0Lh���<�*��4,"�y���'Ii1���-��蚶1�����F���]���I�W�]|E�0�{�dM��ᶡ6�������������~�$d0�����D8W"%b��[�R���3��|�ؽ�IM�6� Ɂ����aۼH�Ze�ؾ#.N�����f�@���r��s�
�hd(����Io�j<���zH֛�z@�ɩ����_�uE*�'�V�ap����h��;�~c�(���!�M)Oi�)gt�]Lxg��	���#��g�0��B��v@*f���0�,  �K���J{9J��p;��ì	�_�y#�@*���~�i]s4���Eh�����z���{��'��ݗ�����J �s�+�����$\sR���*���p������Y�0���d�,>��i����~�ڼ�'��=��0R��1�,��I`'�#f�`��CUj�S^���D�;M$4}���y�<��0�48����L���M�qb�����BJAQ[���a�4T�h@���e����Y嗄�J{��+�i9�%�ǢϺ_R>c�A�$ @�P0A�#�����s���vr6l�HPFP�i�2̸`�@�I:F�-J]-8�^�h�?a1�n�)�fX)
��5�y��UD�t��@< t��e�悙�/��n��i���@����������i��ԡl �?��BZ�mB���v�~xMDے�3|Є��;S���`���	�z>Ø��KK�ٲr�'Y�k�[`!t�ųK�P<��zK��:m㞛�0@���EMN?$����}�A(�V�����F��C�I"���BC{��$R��KQ�$�?��?�N|����xC=���ql���F�]f�tK������ֿE�9ת�Ϝ��T�i[Ռ�����|��٨gU��+��@ZV���Ģ֧�LN�fY��'�sSvmZ�q���Zҍ��!mx�w�!0���3�DGr�(d��(q[��,�ַ�Cd �2%�p�A���\5H���ZY1�l���Xڌ*t�*��;<��SH�j<�+o}���Mk�ە�1�N���xe�G%t�kk"�ՀSr��y�B�kίt�_$��oZ�T���2eG3X)~������84FL�k��o�-��wI5�d2��jB�g� j)����/"�kS�8	�UА�kbZ�K6D�ǏZu�H�\�hc�ɶ�8�p�}��G|)d�t*Ȝ�=q�'�yy�0��t��
�p��*�)A,�E!)�[�w@Bay^����$��we8V����B�\-� r��,!��>cH8M��o�)�*�4���8UJ���"����>���������`*��p��{�n�h]Fg��0T�3d�f[r�*"��.�r_���iF<�̼3����ƆN�p�������N9ݸ��ք�nI�2h����&~7�~�e)Q'�����{�Z�a.J}WʉB9���N�-��v��of��.�\���U6L�=�Y@�7�	杀�s�Uw6-ƽ%�4���@t���� �t���v`����A����h;X� '�,�B�E_���+iC�� Q֖-[�q"���f�w�}7�ꭈ���]zŒ�+
�3�Z0��c�m���)�!�2)jUs�>zu�˴j�f������B��*�'�d��� ���B�n"ɚE�=��ә�/]��c�/��b^#m��<4@Xw����X�,���*E���v¥tՁρ��'��`��e���[�lP�����h�޸� ��6@���qV�KX	j�����p"I����]��oo�9K�n���҇�p�g�r��C sbvG������h� k l�"�J��o����"���z�N1(��g?�g��فo�n钥�Ϙ1���-�Od�@��}�m�N��a�9�DGqgQ{��g8�/q�ೞ�Lt�=��eˠ����y9�H���̝;�Se"���{.� @C���+3���Id�Jh¢/sSv}����8��4��+���� �C�âYn�?��]���X"�$*"�� ��c��At�_;���* �&v*GG��L�P�&Gl�Xad���^����_� ��!C����f���������d`��X�^�#�Iރr {B���7�#m	�Z~�u���(�Ţ�@ =fi"���K����ԔT:� l��_�}���~�#,G@@���`1��*2��5��P _��H U�.p��1DO��'>A31�3v���B\_"���9܏�2��rHY��p9@��\記YAzB[@�]��tNY]��㡝���@��"3$ee�r�p%�D#�L�P�=��,G �����Ѹo���� ��� Z�'�p���>e���.��#���o��wQ?�I��aQ�,�A�(��K������Da�N!k.���������*΄k����Q%�����'��\O�>���4��;DlLD�C�d�PD�����
d���0�E�
Tc* �y#F=LM�^R��K�!t����ߩU^8�_���ԡ����ld;8��\>���%�\�!CX*�����}��%K���mRd�9��) 3�E|�S����v�1��M�N;���c��Vr�UU�q��X,�5���;bW�Ry�GÇ��XĦ��ZY�p��/D�\�n���|�v�,�3X���e¨�,�3�=H�'�fx�,���5D6�mao��F��xa�1�	x�&˜���%U%�@�8� g J����T ��~ɒ%�DnP�)h8�ԝC����TO�>��< � b +��#@�
"
�a!0���`�0��V}z �Tp>K�K�'��e|�녕��(���'��@���_�2;D���_���R�B�B�<����z4ˠn`�f��lS)��^ �x����\���� ə��y��S��0��<��nm#��`�g��r�,[�凫Yjǖ#`GHP.�.fݲ�	��N����-ā+�D��, ?p�a93��s�B$S�/�؆t� o\C4gd��k�Zok��40av�%�y�V�!�l�Lp���P�9��	���'�S�0D��Y��\���7�'(+�D��C&\N߶���YйY�i�$�Ơ��^��e�{Ǉ��$�Ph��b t��:t]]��t�eG�[��ާ�XE_q]$ٲ�g����6�+���>�H����O���d2"ݫ\&,˖/��"����&��>ș���(	Y����I��y�x%۱	pd�W��C�Ůz����f��ZZZ�U\�hغd�H��I����Y�P�*B[;��0�3AR�Ĩ� !��tS�o�ы!�x���YY'M Y�3*SOa��T����5ϰ�\�g%�@Xr�~�_�A���$��`��uG�����>g���*�L0d?�]7�0���`��o��rx��͡T:N;��T"�æt�#�Y���#��K��]�i�0�> [w��e|q�-9" ��p,�?(��^@%O��6���r��cP�h��%p
3v����I�Eڧ�ƀ	?���rn�AxX��R��јͫ|ȵ����8!vLX"$� F,�	�a��sNd97�w[�P¸zܱhi�����0�$�A���=���mu��5�\���!RF�@tJL+1E��/t8	���<W��\=��l2<8�l������C��R"�A5�1���7�ܴq+�{]��j +�D��^��v�A�|-&%S��{i�^�s?{�u�ԒR"%G��GV��Yl*� ��ñ��U.��LGw��;y���`�K"/q��;!�%�j� �=|���`-��6ᆭ�~��`�X1��fN��]�og\=c:� �taǨ n�Gc]L��ٌX:*�?��;CdU6C�u�P���U�r�0�10"#���zv�bօxqL)!Q@'�|"��s�� �@���A�lbׅ$Y�C��9���h��u��h�ȱԶ����p��jK�l+F�T�b1�J��uS]}Ŧ��9��Z�#5�x�J02���1���3�z/��+�T�!2c��U�F��p��X�N��	~H�S�9�1r� �����B$�,۶��dɒs*΄�un�d,�H&�,G�1T��e���,�+��l]W��eDp��	�ʻ[��u�2V,���2��v�J�V��<���s���:��О�1 #h^��Ndv%��ۯ,��)�) a���L0�%R�t����9��葿���珔L�����*��cQuM�z{6Pu�G��z���C(ѓ�_��z��)�Ĕ��L��uc2Dď�U�����aܕ�`�~�w�ل��	�$4ъe���
ڣ8NESFy:�	��H0a˲lii9�� �sЄe�\Ĭ�c�;N���=�~C��
��8.���d�:�fK0����G/`L�WʔN���!j�,��rv�֡i���Rs��<{�ˬ �UO���"4�B����5�j�אَA��ɁT���>���2S»�1�.��:���9��mS7]��[����J�]1�u��^&��&Ǎ�at�QG͢�.?���g<|���t٥Ki����%��5̂�b� <��S]����aѢ@�\E��6+��ܩ/�2(69^pI�7i���l�I�H��1:f	��94 �V�q�����2�z��{���%2�	x
��ߗ��) ,[���6)�(z��ש������ib�U�4ȕ�`�|���.��v:7Tv�Q���\�$SNc����k�ԇW����g¶��pH=Df͘�}�������"v����?�-]s�w�Pu�Jۈ��{��ldQr���I�g>�x�}�Ewu�袋��G}���*r=�c��k,J$�X��\YP��d�:���-s?F�%�q�m�䵰L�0a/�����#����I����t�@'f:��g�l9R��e�축M���qKȂeY�x�p!���B�uM&�u �6�_#��} ��ʕ�Qo'Bf����=�Q,�_i�r&#)����B��v�w�E����g����R���5�G�̚ <�H���{�5��X�%:`�T�x�G_��{tǏ~C�UM����2c̮���6-���L�5)�s�1�ŋ΢Q��y]��6:����Օ�ɠ:R^�#"��lJ�:��[p(��_1������:�LT�U�~�1��YO��@X>}�\,�N��H��8儹��>;�{ ���/^|vESY"w��0{��ݖ� ��;�@��]�{[0�� ��gJ������Jf�1И�V��#��Y@c���Y�0!�	�����~���e����2�DF��ش�t�Q�i���я?���wQ�WQڱ�@�Z9@��z=�϶�]<����(}���c��x<A���~�ӟ�A�=Y��p�CZt�-�y����g* (���
fFy (H�3�~ f����'�}�, ,�$�o1=#Ć��f�2��R��yB:���+V�8g���{��{ʐ�|#�e��[%�/�T�NF��Jv��F*��a
MES�Ҏ��Q �W����Lt$A��N^�������X�Ɯ��}�Di7����lJ���o��1C�l#�d$)Z�rV��fq��$UW5Q�!rU�s:}��̣����j��t���"��ck�{��0�V�����+G9�g�Ad������* ,�vp��������a�f��'�E$	;��q:���H�l��� �ͪ�m2��
�n����Tt�� ��	O&�°��̒�d�w	�ֽ���v�L�C�꥕+_���8Y`% 1�,8�����<��������_C���҅��4t�8:�������(ք���jiJ�{��;� �I���y����$�4�B�
��;m��! ���]�E� ��C��R2��H,ʻ��%ۈP:��6�Mv����7KLK|b��>�zM�x������;Fk�;�d���S�r������W^ynEA��7j_wkM�{��ә���+�k��#t�~� ���5�	��p�Au���/Ȏ�i<� c�x*�dv�:�7TQ�LJ_-���1�c�Ow��|�^x��`��SQ<��a�r�}@�1�2Ps�4��v��C��I���"� ��ҞK�!�b�h���`��b�����qd9�0�8���L����e�BLX|Stv[�g�.e�\	]�5
�lXo,�dS'�Ax��˖-;w��魃id7�l��zk��5)WtxBu�蚯1��M��5���ܱ�L�|�U��a�r�,���o��+�tI�h�.�a������������
u��N������c1*Ή{�巍~P�m�
��Kv/��f6��������X�gY1�OCԂ5)����Nd������M������0_t �2扦��]a����ئ�{���yf:�f��0a=�ד��L�	���g�BW�w |߲e��ms��Bn�	���N��BŰrl@��)4-�A�s�lp�Ż���� ����~4d���ӊ`�r^�����TXm�r��^87{:�w����6�p�	 �~���ֶ���@��ة�8]�gb`��5�6��$"˦X,B���c>��
̖#5�\_�,$G�kC a>L��$yn��qҰ���Vˢ���F�r�9+d��%s<��[����z��dG� ��,Y�+�rQ`�����I�2��\�U�aܷ|���*�[Zo�IuMB��D<E�U���dG���rF2L9��	�e��$UF�4�lBJ8$F�)�>�隱x�рa(�=�~���2U	kʌȈ���#�wf?�	���ʡd*NQ+ʫ9~ҴȴmjVG�M1\^��0_������`��{$���З,�o[#nu�Y�A��+�-^�'Y��%xj8�1(+���[�`Ov�0�o}�^la�Ul��>#	�		��|�6�%׍S�mQ$bR:��^�8���f�u��B�j^y��yWt7�I���ό��"�r= K��VObf�|��ÑL��,�@�� �x��">�qQV^�~������G��xG��>;g���)��m��.^����3g�L��/G|���M[Zo�%:&!cF��H-�`}M��{:9���C*K ��X�1x8�I<DT@e��ȳ�>�ɑ%яhf"����908�(�
�8O O@X���Y�Z7����]���R*N6�$�IɄK��"v��$�	"�!;
	1j&)ׯ���GG��<����;63ʹɧ���{aq�	 �^�&,;x� ��b�Z�[3�
�w7�zup�{�I�`��L�ӎ�d�d" $n��V��Ӧ��CS�΢�j��E�[�|v�T�([v�f���|���g�������I��?��o�C������f���M�G��yG ��4Y���Y:� l��T��)9,p���x�eݳd	�\Yn���͵i?w����1��������Q�|C:9��|"x�Rا	,�Ǳ�',T�	�׳a	`JN
+��4}��.��z0v6 ��� ����Z[_&�H��ɱH�5���SQr�AV���a6��4��5���;��wH�[by�Aٻ��e��LA��_�`c�`߷PފK	��[a�,�>�Uib� ���-XĤ
$�6* ̣M��/X��*�T
kO)j�4���jklNs���U�`󇣨y�Nd�H(�o��,Iؑeq��
 ��aGu� F=l3����^z)��u�]�dO�S�Dx������ ��^�L��^a
d�Cy�+�c/L�+;6k$ϳm��ŋ_0k֬u�i�E8�޺��LO�TrrG $�����9���7��-F	<��p]�Qd��4 I�![@w������h?�F\5�s` �k��H�P�����w�R0:���^��Y�G)J���ݽ�b1?�r�dU��[hŊ��֭.ّ*�.Ǔqf�G~�=a
��.��ϻ�`���X�B��̪ �U��g�@F(��} �K�g�jx	(@X��更����a�ʻXD�ʤ�S`�!>���Ѻ��ɶS4���>�S�}G�1� �xJQ]�pRf-��DK�UWײ��Na[���i�O~�LĂ�q�㫯��������9s氜�裏���!���?�C��ȓ�2������%��ʲ;������������>C���D~�hѢ���-grOo3a�0nn��It���M��x�Lx2���3B �� %F�5��7��'d��p�@�R��5���������>%Oh ��K"��@��������˒D�;�V��$iܞ�����s3E#u����􉏟O7C��%G�)4g�?�|�(���������Je�ʻ�T�	�re#�j�GH�~N8D++�`�>ɏK���m�4��0�a` @�[��6/ۊ���Nx������G"�륆Z�/�O��9��V�����^j�HS<aP4�@N��>S��z1��� ���G�!|o���1c��y���/2�A������П����7�̒����@`
��P�ꃄ�M�I$P�_�XX|Z�C� ���{�e�����"���-Z��� N��z/>L8��s �O��#�|�?|c�#��9�0ȊC p�]5*��[��Q놁q�:�(:묳x1��s��N6�mI�%+\p.v�����7�N�����:=����F�l�̙{�n���xo�^}i}�c��4���(�d�s��t���e�roO�L�����!�����E.����Y�pL�9����|W�����;����;��Z3��E�E���g>��O���sB�P�+_�_���DnE�]�x>�|ұd��J�ko��g�}�&�=�jFS*aR4VO�
R��sv�0������a	�����?�����3����d�©��������'^ G`ta`
�駟�~l
&,a�����*�u���E��p�������.���-J) �p�*
��˖�	E<"v-��1��<���]�7��Q�b�|������x���l�=�k.�M��\0�O<��xE/��B�
]u�Ulp_���������׼�y�vut��W�ڶ�@sN=�.��T��W^�Dg�u)�kMYu���r��� M����^-�(�����s�����Lh���\c _�/k �K��cy�r�+.3���}5�c8���� {����L��,l 8�;���;n%�레�K�z!���㑏����7�u��]���i��#(��)��D5{^�}*�YL��3 m���C��R�8�́�b��~.�
�|��\�8F�_    IDAT,��<��.B�d����?:�.A�����cG�O�m۾kѢE_�(O9w����kni��T��g1���/Pm]�|������Bb�͊sM �����(�P�d���=v^�f}�H�y晬A��/}�G(� c��C�\�&�r$װ��E�o:�����詧�JӦ��o|s�3~z�����ͣT���	?�
�W`���79����Qc������k�>��+K9V��a@v�eÅk��8�xa}1�3�%E��tr�i9@8��JU�-^|}��'RWw;-�j=���4z��w��4}�!�(Faf重b"�%�����u���>��>�Cd�������±���+H��ԧ�3H�
 �z����(�ɕ�<�(.�!�\lf��������g�毮����}ϙ?s��ͷEz�L�i~�F���g�m�z��'�̎�_q�nZ�P���#`D��3k�,�X 3�%�~�1��7�J��r
_���cP���Q�!1J�%�a3?8���*<iX�����+_Fo��53i�U���L�Wm���9�M 8J
��(F���~���AKB�B .��#����9����b��$1��Co)=����	0�Y��~��[(�襆FE�_�Y:�#�Gt��W�SO�Ұa{З._D�L��'�1���Xq���L;���J���z��N:�N:�L��K/�Dw�qmذ�/^̑7�x#/�8�/q��%��AV=��2�H_��@��������~0H��tJVṑ����._1��ɓ�Ʀy�#&ͻx������${�q�]e��	��=�^~�Ez��g	���� ¸A	'��1�'`(h7�
��2�
`��a��g�i����aA�q<>ñ-Z��� �qMLAp���>�������t啋�����A�^��&Mއ�{�u��GϦD2Fi7J�YEdD��9gp��q!���Ǿ�,  �曯����	�vwSuU�/9�N��<K����7��'��iͿ�2�c�=��7ͬ��N��㽝��C�����А�v/^������s��	'��}��?�}���e���׿��H��={�l:��=��;^� 	Y���υ܀������G�����M]��
Ѝؑ_/Z���Lx�s/�6r�[�ե�3"xISt�!G�	'|�{��f�2]dK�%��������L��w=='�PBBB "Hii�@��҂!�8���w����f�$� ���)�؝QQ�+�9m������OǓĐ'�u�u��������_�~����?DfI'Wp.L�����Z���p�҆��68���"|���P��r̄�6\�n����^��]{�n���q�����[�ՕU��R/��1��� L����,C}��%�9�t�}�*�rjk-k��߫/:5�y��g5��V�Ԫ[n�Co=��`�V��4�<M%��7��d�~����[�DE��6��;묳�S�����'�ֹ�q��8�Xm�|7������8�b�s-�n��N}���3�ל�r7o
�S�V+�T��;�ν���L�8���=fӚ�z:�F.: |��O�y�[?��g�a��s��7AB��:�!�r!�)��@]��Þ�|�K_
�{��;<��0e p^N'�fr8�c�%�s1~�bHV��ٮ�������Z��I����ڔϕ�nMY�w�r���%Ӥ �f�$O~G�?�����k[�e+���^j�&}����E���Ƥr��^zq�~�����7M��_?��_���l0fHS���A�!l��	����)G�ڈ#�y�����?�A0G��7q�y���d			"�t YH#�P���+w�h�r79`���4L��JWM�SO�}�]7�r�)�WE��o9j�����Ӽu�1�1�2�������^�Z*�IPI� ��TX;�� k5�5�����Yp�q@�^y��9���<,+戾��t�؎5��Љ1�=!$-�}�7YU�	�Sz�!l	�U���P�{�K��1�C��ɪTM)�	��4y�t5n���!~m��P��FᕫW�Ա�CMMe�}��5mƹJ���Jjn��[Kڴ9�|>�Lj��R�{�q���tD/%���1�Ad�=��}�X�17`�%�!�c��v�i�q���6��"�O�+����X�ҥ�}>8���Y�|ꩧ�y�ۄ��L���wr��Q��lZ����?��,"	^�a���ks�F}���U[#��W�X\p�/�a�e�sh �EP� :��dђt�+B�q�� 1��s���}��� �j�☳(�����\k���y��[3*��)��kX�H�������ھ����&>��*T�԰W	����vH�	0��s���@�ZHh̨V]u��z׻NR6[V:ԆH�\kTwgM�T����*�Jg*a�Ѱyp*�+~��<�i��aj�[�xm9A�7���G bS�N 68;�u�ĉ/���f�,0	��h�+�=�F�tWOwg2٧�y���0~Ӗ�����yՂ���I�#�Lވ��:u�8t����3*vcG��h,����߀'�^<������9��H?�&��q�{�F�5? 3�����/� ��a���X�`SvP��s�)�8kz��O�k���BO��P�2���k�(E�rج$N��K.�l��UO���x���P;C�/��C=��m�n7ftV�U��[�m�*U���ǝ�7��r� ���BoAz�I�,[�kD0�K���#����B�0���ի��;��N���I<'	Q����w`��8��`����ӟ�e���V�@��s�D�Z%c�s�����xío�i���|׉�d-I-��d���Stҩ'襥��r�������z��:i2:	���Fh/����C��6`�>���SO���]�Vs��	6c��m|7(�F��6M&�N���gU��:gRd�P!��>U�V�V�as�ƍW6C�r�@�Ƽ��kH�%+i���Tʥ�%ns�fʪVzTKBrjjl����Xe�#U-g��ܤ���`��ը�V�K�
[454(�ӼP 8�$���2�!V�����,=a�u�5��H����P�j,�v���k+v�&Rۃ�@���.����j�J)˯͙3gp����_^�pT�<�;ߝhmjU�3�7����2���5��g�5k��ES�ދ 錗f� "��I�-i��	=���3_(ڇf��@TT"`��k,���7�d ��q�۵t�":+��m-( )_`Ś��F���QBS���QGMP:�[����~!�PS�Z1�KOH�FU�Ez�N������6��Qo����ViPKK�����j���z�p>` ;��9	V�z��a��s��F[�3�ӎ�]̙�� v��6mڴ�z&��2�{�F6��ɢ�j���}Y�qސ�k�H���ܹs?4�E��ћ6,l��6)�I&��/Sa��u�X������MZ�|e�`�m:�"�N�0��d�j��x�t1�`r�Y�pZ{?h6�f�-溸� �����v����^\[��|O=�;Ö0�P*�6B�Wo��a[���
A���Pt�^����$`^�v�>���T쪅H���4jX�O�Jgq�Q$�Qg��B�:�ڢR� %;��)U*�@��G# ��w0�����vK�-���~�^"�LxhBÆ�]w��#��v];��@���8���xa���MM ��G[Q�"HP @�v���Lx�A���ͫ4to?���A����2h��*��:�Lw�[C��@��8:�Tm^���/t��? ��cE=���P%��% ��DG`~`9�&ta��"��7�!8�=x��xƌ5�(�R&�m���eU,oWKKB�JR�}~�>��g�eK�������Sg��!~���P�Q�+����ROU�nӬ+/�9�P�,�*�H�FU����u�R���������p?Ha_(>0Z�����?���%�)�6u�z�Hڊx^�s/g�b����Ŧ��z�OT��8�_	_m��QZ�M�6q�������	£6�Z�Z�91�N$�@��F1���+ۘљg���?!�V� 1�s99k�g9�ҀNq&�t �������\G�������;��@��a�$k��w0�2ib
z�ڵe�
e(�פ�/n��ݤ��ʵ�  L���(C�A��C���%�	c��֥�6��;ޫ����/D���`utI��P�I�r���l�`Xg�;|*.��5~3���RO|3���0��~z��:m��!8�� ��?f��W↹ ��~��6 �	��b� ��x�z�Q@�����Y�R�>��J�mI�=eU�5�(W�Ѱ�vM�0Qd�'L� G~��� a�t����g{@�(qu&�
"h�9;��N:�t���(�	;N8~}�a�U*t���򸎞p�N<����Vuu�fUQ^p�*�*ײ�
E|�N�g̑m7��=V5pI� �b��������'t睳t�{NUcSJ=���,ڬ<�k�t�jh�Z5�T�1D �{��f�@�d�x�3�Y5ϛ7/�%����e25�1U0�!|��<G? �|G�	��s8߬����^�S$������O?z��7 VΟ�H�Ά����	�E�a(��÷�'���cJ��@g)��vT#XG8�e1�D@�|�^�z�i�:���	�Q�o�p젣��|�>��U�nҥSߩ�o�'w,]�U�\t��y�8U��as�	1�}4Ǉn��K� �d�KZ��Q���WB��E�X�����O=�mۓ��#Җ��f%�ٰ�'�!2��'���C�U<d�3w�4���js]	���fe������������q�iq���^�Y���+l�؀c�2�5��+�L��a����$%��b���d��锺J��nKSk�xd�@�`��~m����(��L�^��pq�����ý\�Ӷ�s�m���r;8F�U��z���ߵj9�[>�����o~���8L�����qoђ%�4����;�r�A5���h��{A�%�s�9^5oH���r�r-|l�r���f�ϸ��@���������G��YW�_o}�۔���Ɔa�r�y
q�3�	c�c ���A�^ۡ�����&�l�^��`K���ڮ��u|/�
�����*��s eL|o_�K#ĵ���e��|�I�jI�M��娘��R��j�.0�t��i�5���BZ�YPt֬�5�^�g;��m֖|g��� 3���`Ψ	�^-���S�W�Я�S5������'u��oՒ�k4y�U*{A�-ﳚ:�
u�ذ�V�N���e�탩>t��Ua�'L�Rʫ����o��)S���C�S����>����;5~�DQ��'_P6S�=&���B&,)��e0����j�ؗ?���x�k 2��:'�6f��zTŰ��ͦN������Lc&<w�����>$klX�c�$!jDG�Sź�y�j-w6��^P���ef�d�8Y�%����~I�Ҡ]�j5d�}|��ziɯuđc�����z�����+4c�u���ܮD�[��2�2����U�wr(cn_�ܡ{�	$����+ֿ�+���pJK����Y���i��>��Y�>������}�k?Ѩ�o�-~��;A������j� L6m}g�N�c����v�κ��{�|?��jb��cL�ܸM�f���͛w��g�mX�������
q��Aة�����}9�x��������{�Ś�O��������#ںu�f�:O7�0]�����3oԶ��pk�'LL�)�4~JgJa�!ޗow���^{��Y�A}D=]���V�w�O�M?O�B�~������K�])}�c���'ջ�H�B9��-��Y�9
�p�R�o� ��c9D�^��b��A�D�7�HV�fD������AQ;�ڏ�i�5ZK='����� �j�7��� �|�����UԦ�ل���ZY��=���}DUg�}�F�N���G+��t�����=�a�Tk)M�	O�4U����ne��yod0t���0^�|��?����jn���s�Ռ+�W�ԣj%�_ܨ_�b�Ǝ;A#F�JYJ�YU�4S`��r=.��)vְ����4����d���w�}�*w�-o��养ao�=� K�}l+��聾�0Q�'_X���_�����8�Q�G��jQ��ujj��UW\�amݒ	?�Z˾]���
5��-1�;T��OC��Ax��5Z������̪���1W.v��+��ھ���N��ܤ(�re�)�lP�R
;k�����p���S��?N�ʌ�k����o@�}��ڊ�	'2G$E��]Oe�A��(	��q����c���	B����T�յQ���RIjWt���]/<�^s�}Z�0�j�b b@�>�O��q��Z��S!�|H{(�Ϣ����Z�i��.��.�{�ijlH�ɫU2l���SU���^�;���K�P}#�L�Qq��6�U�>X <w���M&�;��S؄w&q@�^�r\_m�?8�b�����*�B�����+�iR:9J��Sc�p�j�&߽�iS��رG���C�O�@=m9�UkW�GV��!ky0�Imm%TV��h�v54���o?M�����&�"��ެ�z</!a����Ef�3G`t�6�[����&��:l_
�6�P��������c����'�DU�D2�B��5�kUw�08�F�*I��Y��H�bHN���X/6=d�ؗox���V�����];b��Ez��G�(ה�+9�J��	Gf\*Ѣ���&s�Z�[U��C"V!_	)�6E���PwQ�cn_DZ�c��L&��3g�����}Q{y���RQ�QwL����C<���ŀ��.��xa�I9lj��m�`�d�lZ_�(4Q��0��,���5hh�	Ke%�)M�6Kcǎ|� \���9b_�١{�{	�/[]�rc��Z���
ʦ��64��O�y�pr�a�XcsV�JU�JZ�dF���1~86�ٲ�������5@��s�̹aPA�^Em��ƞ�I�L2�L��</�&5TC� �ɐ�P��o�+�;x�I!s�d��x@~;��Kg�8l�b����f�~�xPU��������[�D8K��̏�C[7n���w����jZ�jc�u�$`U��-;c�<����b�	�\{���^�������*��C�Ր��!#JE�4�T-ըc�9Aox�[�/���w���Q�=��!i�#�N��3ژ�$V�)��u���%��9B��;l�����z�	�wY��Xs�1���Y�={��&MZ�'�m��	7���Q��>z@�vR�Г`��T�j�j��/�Ԙm
v(�BH��3��������s���:Β3�v�˲c����]?���7[-M�ri_���/&�eIԣ��uИѪ�s!d-�j�ꕝ��;U.7���3�1���)��פq�C�{2��ݟ$�w ���Z��Q%*y�SE���t�{�PKK*�(���`޺5����a'�R1���ȐmZS1wg�1��/~1��Lc�5���ט��Ǽ�{�����=�'��=�s^9������9(F��l^op  ��ٳg�8� <fÆ��ʹI�b.TQ��O�TT��U0ឞ|p�F��|�^.!I�����`r�9��zI��d��C���Y�X��ls���F]uլ���	����Z�ڇ�4rTZ��F�#_]Z����}D[�$U�5�k��ڛ�\��1�����O%�`fL��l�j�_����˦{t���5u��*;B��D�U�JV��m�-*����ԔN�����ZNJ��u�� ���BJR�<x�8��} n���w�뚓K�� �WٜK�`�Sٍ�c �[:ǳ�cP�R��R��x��M�8��=y�d��|����S�7M�6�m8Ԏ�]Y���*�dGӱ��%U��=q���t�P*�S�3f��k    IDAT�6iX�,y���Ջ\���Z���g͚����3`�����n��'���I��q�^wp��wvj�҂.��fuw��Zk
*�	��P:��VJ[ޓ7t��	�q�=�ϪV:�ؘ׽snԥ��T2Q��=�\������c4|䡡VwSӨ����H��|�+�O�	�1��l�%m����:+lr>XCUF���!���� (�&x.�p�����JYj��fJ��ZĤ_���a�fV�v�̘�+�J%�L>����4� <f���M��IM쬑/&�А���V5�4��'��N� �@~��0A�ri��v �E�@�)=���?��E,%8�=,���6wxGf3c�-���؛8b�QJ)ו�,{��t��g��NVk�0-[ܩ�fݦM��� \�ԩ�â�y�:d���+C��	�W�Y���>��6���{�����V�����>���UwwR���7:�ȉ�犪���S2I�r J`U��Ļ�Pj���
PdU�R��}�[21������� �ls��U`|�ƦL�(\�l����2����N�j�
?y����t��n�Y�	{�mG�oZ3���cgQʒ퍊ł�M�)��]��rZ�	S�޻�� W;�EP|:�DA�z�O>�d d�f��jh��m2�T��v���W^yE=@<�x��� kI�[���KK���Ԣ���7:���Ӣ�o��iׅz�;@xGQ�T�h�8�����K:wH���K�X�D�y���m5"������s�Yڶe���S����ZZ�wާ716�0cd��u�H�����  l����/�2�l�.��5��~0�x ��am�q~���N��g� �"�`��^���f�@�� ��`���7���~����^�ʃ>��Ae��m��7�t�H(IC�I��]��&�]�>G�-[��q�lH��C`T8�cMf�(l�6�c��^����4/�v�P��P��[��V�F���"Dvr�:ur�vI�`}fI�ۺ4w��Z��Eez������3V[�t��SU(4�"�	�{�	_��L8קþώo���=q���?J`o
��¼]0�a�6iԨ�n��Z]p��ܾ]w�u���!�����Ə���C��r����|T�/�~������3���g�s�'?�I��:ʁ�������^q-r�6N9��ٟ�Y���e˖ ���`��s��ζiv�`�
̨�<�LX�C�= �H$���'>q�����7to ��ܦbG^�v�ο��=f�^��"�Z����P2�A(�Lh�p1`�!��ݖ���ǵл���`� ��t����p����aՠe{CM6�+��<��CT�@ǖ-���}J���Ot��-z��������/,ѕ�nPG7 gBhM��p/��,�K����N�?E���m��u����Z�r�.�B ᖖ�f���f̸@=]ݺ�������:\7}�M:�4u�t+�a�	".=����6�\����
@���؟P@�`[2�U�\o�����??`&-�9:�@�U�#��3��6p�o~���S/�+'��'|��[���8?�u㉙lJM�-*l���<C���4����Z�z�:;��	@"0���y{Z�����#
+��1� .����f�N�%aI��,0i>f�ZL3g���,�ӯZP��Mw�}�zz6h����ʫ.R���z�՚:�usD�pR�DF��my�8%SDGTT��ل�h���x�D䭵c�ks;gm�w*�\d;6�Hj�kCk+W���gU
ݡ��=��W��|���o���-�'���l��#�Go�t���J�e��2��0vWp��N~��O"Q�!e�(+p
��7�b���WVӧ�v�N>��p� dmN�M�.���:̥�.~�r��`�t0�(���N��<o޼[�&<b������]ԝ�.�l�|���/~���\�� ��h��.�(<���Tl@����~W��կ�0m.0pp/<�쪊M����Z�e�8�aq��;k8��w^�d���o_�!�������MU�	�\֡)�?���&U�TQK�p�@��{��a�)6�;J��1�����"�����|ò��=��(�L�1�Z�?I� �l�r=���Ky��U���/{�e)QYL�w/lҢ7�u��S۰����Cj��ke%��Q'P�	������}V˄��{K��r=�~�<s�k��N�0hB�p�a�4�3�5p��
��/|�g�������o;���
sD*���}��w렂0!jlX�`��'�+EU�5�~̡�����m���_�,DX�,&L��g�5�uv	�H�8r��^�9���P}��![&	���/gZ��bc|l�Ahl���}��f�;c����9"��L����ש��M+�nׅB�E55�L�P;3J*�[O�7����ncfj�J;�vV����WVT|�跗S�����u�ܟ&�P[^��KC5�	ko��=KS���&Xn�r�mڶ������{�3�bK�L��(/W��W׀����0����-�?�;wn����W�vj'� e~c&��=���e�L�6-��f��0�AI���9��7�������L��G[X�s'�Kj�Z9�J}y�A�����ױ��-�Z��;Q3g^��|�b�k�7�~����+* ᥮�6tA�����da�x>R;� ��.�(�{�����6D� 8K^ ,!��$��}�{Ò;���	R�J�Q6-�z��mXV�|I+�n��om��S/e��׉�6u�ƍ=��9� ؄�|�q��+L7���)F�x����7d��p:�$���;���>]��i?���I�$$kZ�j�>:_���F���_���91���
#�+�ʹG�\���L�;bya���as&,��/�g��v�K.�$��(�M��ډ'���ް�x�A� T�;�j�S܇U;�8�29�����=�d�9�;_��v}f���D� |��'��ߣ��ڼu�J�r�	�����j�%9N?��p��A�'M�:Jx�w8����s��9�ӷC3���p�eP��=�RHX>x�/���� ����3�UWG��Ŝ��)<]P*1LK��UCK[HJ񌡨�� �
	��W˄��m6�2���"!N��>�]6Vf�S���
����r�I�^d����	>Ԗ�_�k���{X�BV�ZE�N����o�ӓ+��Cޠ�O����R��U�Pϐ��V�Ř����g�������k � I�*��m�g>��w��L�iچ)@uL���� m̞�1��8D$q˽��1��=��s۠�-�^��ݖ)����E]�����Z�zE0G ¼�����$��!cǍ3T��a�,3(t����2�����-\^�C����͂����aN�EQ/��H���PH$��A�Q�@TG�
�j��ɢ*�h�:Τ��I4�^��L�]~����'���z�:Q%����8+XA`
r.���1+����P�'	�A��%+^�#_���ڕĴPٮD�:UjUe����:b�jic�܆����)��T��ѕӜ��(+��0q�_}��!B��9��SO� �c�k��� p�;S�8c"�i�c��ۨ��<�Wp����q��3��
�ͪ�w��={�-�
�0�Q�V-l�&aFx?J�_>C�-��~���X��P@x�ĉ !a�Ȅ4�S��8?��9����`� ���Z�[Y#P/�]t�!qQq�Hl�@�uf\Q�RԢſז���I���H
xHM�����J� \Ӕ�3��Ã �������~����]B�V>V4f��ӡ�(7!���q��4����ڐ�Axպ���IU�傚�j��u'X�Y�L�&L���*���9�&\VR�>s ����ς��9⪫�
�"A�0����>�g�� <s\�0O=���Kd[3`��ò��y�
@�{::\���b�zI�O�}�݃�#7�\0J���{:��ԪCF����J��.���.؄q��@v��4��q{����YN����l%�&�%�� Ll<�=�%��
�հ���̆�X�����|n�~����ٱ-���
��4;,zi�jlł�!U7GL���^N+E��^�1'-O��񋱩Þ\;�,[�}���^ �d���V�3^S����l�X�f�}d��]R[S�ڇ�Ԑ�&��Ҫ�����>H�}�:�����@��WQ��	��:v��7懛o�9���8��l�Lw����50���
��|�+�r�����(!�S��p9n;4�`�&�����L�"�&�V�~�{�yP�	S�}����O���H�5F��ݺ��[B����%55�v��O%��a�6Nl,��=��H������;��܀V�		AЀ5�<0;��0d�H�6Q~c�L���jG�T
�Aw�>���*�rJe�J%�ܯW�{�B��I�T�M��d�: �y�;�#����8j3[�G3#?�o���f�^p�|lj�o��6d�(0;��"��0#��]���-�J���%����0bs�����Ǳ؁h��a�~|��!�����'c�o�e�p��WHV�nw�3���{�zEc�eD[�N$`~���s8�=��8}�m�A8��Ǟ�O�?/�}̠�7���dM+V���?�\G�=x����<]|񟅚�L�
��R�vmڜS��c�=��R�=�ݳì�L�����7����I�/D"Z��<���{�a���+��2� �I���	�x���L���yLÜ�aA8�o,��p:�~��{��Ƞ�1��Ft�_���v2���������N:F���i�˛T��sw�iϧ�;�&�'8��d b�AS�>Oh���_l�a �����*)q4��>8�x�Ax�ῨJu�F�H�o8D6����Y%z�5e�5�盂3���$l�퍨'����%�`�������	I�\�;u9xI'��~����'��<ϓ؃� ��������!;?׬����:l��\e�fE�wo�j��~��ab��z��������4էhl#7�������0�8��Jn�{B�
.vj���2�ǲ1X��v�ڔ��ξ��&������^���g��n��ݯ�]�A8����ݥ�l�M7O�ԩTQc�5dҊU�U(��N��(-u�&����=F�.�>�\sM`�8�*�[�2�����o�'Vӄ��^����&�6K �=��9��Y�C���>�{s�p*��ڽ��{Ӡ��ȭ�6�t���ܐ��O��:����i�Q�!��~�֯����^BG~tfANU�0�J�޿���&����� �����n#�'��3��L?!z ��z����|�T��%U��o���ƌi�{.<C�-���V,�Ԍ�7��3�J�Y� �鐬1n�X�ӕ`SN�2�k�>sG/H8���qW}�9^5�@h6䕀��`&�I�Ak��{�fñ��@36+<4?�7@���i{2h�1ӴYē�>���ǌ���d�x�?Ã����m��=��$���f� �^_���&O|'�� �qj��L�tr?ڱ���឴��oF��gE�1l`������"�?׫�6� �Y2�e+Vh��_P>ץ���u��v��J%kھ�����J=��M8���%�J7dU,u�S�EdU}{4�.ή�����#��E88
���г����c.��� �ؓ�+�>���w��x����&L;�+˲w�� �9s�|h�A�mÊ����I�R>�Ne'�	�x��B�U+VkѢ�B�bVeA����d<� )��x;��^f�)��{�qR�@h3#�|�|�p���\G��N�Ɋ��-�}�Mںm�.��}�P*����AS'_�Rq��զ�-'�5u��^.�F��pn%l�֎R@�xbz¡L�rI��X�<�e�cv��;E܊�l��f�?�gGGxBs-��خ��������0:�ȸ�eO ���cFƳc`5�5Hr//�<.��v���\�UV�0��0�Y&6�+��9�g3٘�ǀ��C�����y�N(B&1��qR�MQVj;Sd|O]��c��(�X	����7�Y+���.ї��E康����;��5����ݟ�>����6���;u�o�鰠.W�\K)Q��Q��`�a�q�	s����� D�^�+p��j�z�������I#��3���๏A�d�c��ް���|�+�1�|Md��j �{�w�AxĖ�G�J'���)jGx����z���j��	ڴiK��X�[��n�@a��	@�{l+[3{�mz�'OA��9္1Q<�< "�)N=��}���i��c�|�����sp���?������߭�{�3K��U����9������ՠ�U��kRO@�(^@�l�p�h�P�|>������sO��0P<)~����;6�&���`�b��1�`�2-	�=/���6��|h�%��Y%�4�q�������+f�1��;���.blvn6�d�-�U�Q۞m���� ����l�1�s�e+�X�Ǭ�J�כ��m{��?~���to�0�{i�b=����J�iB�c�.��L�x�+}����<\��>W�&�j-�r%/��Jg�D��)��i;~�O}�S�= {�>x@������n<_p�"#c��Am��q�U�My�����}�k}�����d20��	صaarۦ��!j՞��U����9g�+쬁p0�tҚ� ��a9F� F���G��أ� ��3L�a ��uυ��	�e��}ܽS&�H�Еל{n����<8�?q�N9��\�E�ϸ^]]��R�0�z����`U��8ᘭ�^�!����><�]��s��ؽ�I΋Ɔk扣�`�g![��#�0}˃ev��1��ywț��0 t*Ê�u=|-�=<�hǸ'�N��`r�ެrP4g<�Q{�N�dblfMi��oȄ���p<�|�mA���@l;d��o��(װra;|	y1��o@�,�y�6u��ܗ��/m�r���ݦ]�*l��6���KȌ�D_9��pQr���h�s���^5�AZ�)�	/]�D_y��ڼq�:�A��1K_r��nަ믿M�^ت<R��:��	jjlS��W-ݣb1��T�T�;�c�W���r3�3�hcҀ���`EO�\ܝ��=8�Y!#gV|�Ƶ�
�W�}������J�8��MSƠ}�8��6MjimJ��A=�l6�|�G�R^��mz�����x>�T��0����[�D��v
�U0�04��ٌ�k�[x+^��`�;�J����V-Z�s��-#���V�;�`-]�AS�_��δ*U��l�Y�t%d�%zkg�� ��b��&K&�MۘD '��53a\����X�Vf"�6@@��&#�8�}l�o�c�e@��� �k1<���J�����asO�E��,y�|��2�20�7?���L��9^�܋PĘ���'�0�xc��!��u��3q�iE;��ל�In`c�"s+2���Y�Z�f�~�����O����˸�Lm�9!� x  &;r����f���`O�#<�c��2`�{�����{�a��J�+���/�1mݼY�����g���g���C�7��S��TÆ�;�Oo{L�W�T�+�P�,YI�o�p��#���{�+f�?Bvf�V&��.�@lvd��EE5�-�I(`wG��G3o�s3�W��
3����aЙ0�a����*I�9loT��U͔�ΦT.��\*�
��&f��P��섁��!����N,x��`�R�����6U�.>3���F3�@��9o1ס��Y��˺⪋5��B��U��1�P��ZkP��P�rf�m9�
gP�>�cS/����D����xU1���ٖeM��FN0 �6@��D�0�,E �AD�p�m�n��&�FG���w�sv�= 	���� ���$���0(�e��;�0��m����?rR    IDAT� �.5�$@6�H�#�8����D��y�| 2���(@�〓MA�=��g,�8�������_d�,Q���x��w�Mڏ�b����}u�
�!}8��2Gބf��b��ܠD+�FI ��I3n�r��(e���嘕;�2xG�p1���|}��|ɲ���Ǿ������G?6C�/;7���������Rg������c���X�E�=�JT����:���y睁�!8"���0����u�Y�>�!3�nPzȜ1땵��e�x���/��(���J���;w��wܚ=��.�7"Dm�5ZK=')QM��= L	�r�j*��s��t���C�����W���IOL�����}�{�+
�Qs}MlɽA�>���x���0�W����t�k�J�lo���.�x�&L�d��&�t2!�=~�{�K��#a�01� L@��pfr1i�����a�ʀ�=��P���z@���I���	���c�� l6��� Y �s̑h���1 �`E�\�5v(a@�~�=?����o�&�p��$�� 5�gs��0`À KD����r$%� ��XI�=�N����
��K{9ӌ��� "
�����;mQ�\K���w��><��slR���{������	#o���j�%��! >���ڦ������ %B�b��W�����0��	�^�F=�9U��P��;��%�OWc6
�,}iS����o9N��c�N��L֓z�+��z�I �E��<�9�E���>��I�.�߻����~;�/$��܏�?��>�����tz���8�L������}�'+QM�)��� ��Hk3/�c��߱���	 <ӶI����&<Px�[��%)٥C�t������s�\�~��m*�S�8Κt�%S�Ru��;�^F�O�τ��g�2alo�\��Ť�@���yLT&�w ,��e��4|�? �hh� �0T 9�,�̓���n���И��;u}W��r��Afk<&L;�:�-}x +,f<@啓��PZV�6#01Q��s�o�t9x@(7�%���\�yȁ������� ������hh��=q3}����N����ʂsQ��$����F�|�c���W�[���{�3s���y���<�N��������Z�2��� "]�s�ua5�ɒ�ߣ��1��Z�f��ŴZ�G���$��)�TO�g�#Ko��1�)+��aj����x�m������[1 ��}����������9��`mM����- ��=��5�����@U�*=��ڤ�LM-�xZ7��Ѻ�=��޿UWGU�23�P�d��u���J&�}��uڶ�6j�E��<�}g�0������1�cخ�� Y���f�_& ��x���ȅ{���]Lfl���
R��"��59�`E�����1{uH�'6���)}`"��@�z��cF�@?m�� �d�� ��}z�8����N
Ϡ��"`�N� ��?�����x��ov~�^0_�L O�0p���C� 6ރK�"G���PJ���D����w���|'�ŃLQ�(&@�U�G���x������A��B��Y�)�}r�(VS<F�����A��3�/_@�1�R��w�:�4���Q����˵�2�[�U��������>���t�Wʴ�Ǥ�v���-�ܰ"�jثgcW��A>^M�'�ƠD"��x���{��?�=}x�������7�o|yA[���;c��t=: ���K�8|� eM��������G{���L���e��FtC�ح���GZ�jE �r�#T�K&��Ғujn�\��i*ժ�L�,LB�t���m�"G��
/ �2��ق�2Y��a��b�9
 `��Ra;aW�B~LP��L@�8�Cl�+���x �XI�T /�`�8�X"�	@�vp-  �rm��.�o�\ c p�]�`6�➀�}(���>� O��p-��<�L
�8�@�D! s�N����(-��= |��ʓ�Se�/rfL�f�N}��<���Q<�����E?�/Ǒ?�@��q�, �ǽ�@�PĘE����ȇ{�V�y()�j��1���x�L8U��W�s=�J����4���?�!�)�F56��ط���y} a�aja��w�.#[V�����$=�-�=���������|��0�o����W �9b@�p̄-�X(ql�;��`�'��.�53��¬���M�Z����,VO��`#.�XK�VmU2ݢd�Q=łҙ������:z^^R�+�/��b"���y�g��� jdò�A�#��a1�3a�,���d�������^v�"����y�,���4��1�Ñ6�7� ��`Ұl��؃]� F&|O;x>��P"+'� Z��A>�>0=;!�5�{1�A��N��L������	
��<��� ��1�hE�;�g�F��=�����M ��G~8�������v:���
�˸�Ǭ���V,���&���7a���٫f©������W��^SK�Q���U5f����c����C_�lC����+W��)rʦ�;~���66��fKc��{��,����8a[q�����nG����>���'��<ۥc.b�;a�	;��>Y�(�X��,�=i�@�Q��9��5[l�B�U����K�
�'S�+�)6m�-J(�|�T���C� �ђ�/M���T���d��H��l��fb���m�LjX8���o�0N�Cc�����M�q�	� ���
L`'4�&�X�k���8 N� R�t����㏶�0a��&;���P�PnY�6Y�{� p�M�<��w���:~����y> �G�0\��=`�0x�J�N>��c<����L �D��6�˱�$ Y E�B�M��6�/���N�y������$��߀=�����3pl"_��&.�g�=9�ӤdwsowLx��EZ��/�g[U�[ڔ�^�D"��l���V+��c�S&۬D�ݐɈ�nM�R�~
�a��g�8<�]�a ��@H����ڑL&�}���_�'g��5Llnp�t��}a�@�N[� c��Db��B���*�.���׆�W.�`�-R�M�>�LI��
�dB	�K/��	&*��Q�x ��0&'툵:@����6:6�D�c@�L�
83��d� u{G0��� �mj�m��^  �( � m����Y���B��m��eN;`��
����W#V�<`�9,�9F���=����8���;# �6���,w�#'�8������w`�7� � �ڶh34���_�k@���1����]�lA�]L'� xw��w�8oLP����L�h2�{s���=a�ƴ�-�w�wC_ c��M�3C�v혫i��z�G��Y
~��ڪa�KJJ��J%[՝��w�Kc��J-��
�j,��|h?�/+{���x��Zy��Y��g��a_o"��&�zd�Θ�>��^^�Z��it 3aw¬�,ƃ��owfwygߛ}9 ���Rʒ6��h_��Ɔ���-jmI����ư���Et�-��'�T��Q�]M�K/	f�x�v��ba�LL �� ��9*�la4�0,�kP,�c��!�����9:"L��ɲ���.C����� �a��	 A����j�e�Ov�q-��y�U����jh&ǵ�����h�8�u���9�	���̑��> {�Vڂ����v����z�'�B��.�ȹ��YA 3'��S��>��!|���Uy�p�'�w��5��
�}��(+l���A{h�c����Q&N�F1V��`�׮���#��\�*QN*�����/һ�}�ʤ���%57�M[�U��A�0�*0ߔ*�Bؙ�J��V�N$���V��_&>�3G0c�F�h�O�7q���}ʉ�����M8�>�Z+'H[����D^�t"�	aa�6w��Zd��A,6Q�K	w>v8q��߶+٫
��5kV_��_D����R:��a*W�����M�^�Ӫ���K$5u��!YO0[��j$�ι�3 s�D9�1���Q0#'� 8N&�3z8Ppvru(��ISbr��F������@�k�T�}�г�Ӗw��A�w�o�D����>�
��(�X����l�ٽ��x2�o+����J7^aœ<fJÞ��<1��m�W��4��� ��noq���w'�px�ɔ/["�Ւ��N͞}�f�|w����0L�B�::ڴ���̳��z�I�럶ܿm�M�(J��Ϗ�W�摝�~_~W1�M\�E�<_8���=�ұ�7[��7	QTs����W
$k$ʥ��eBD�!c{h��D��~��,�����w�b���$/ `qzk��⥃Y@�]{�}!j��j%�[����[��z����Mo�|��߽�^׾�c��ȆR�,���:uZ��T7��?;���+�y�Xi��/��������7��A.�,��c�B^^��)�tt ���q�Iag�.�R/+�|1 �n����w�;c.���o+���p�T�190��0�K,�e߳���e�6�N�1���_�|��+�݁���k���/H�����{�L͸�\%Sm�Э��vc�KG�=Q�v���X.)��(A��2���!��7��x|���v�ج�I��q��oכ���c"bR�Xi�!?�Ǧ3f�i�`\I�Rߜ7o�5Nػ-7�;��\����p�݉������f� �M1S�Ϗ'M�<��3 ���ۖc���`iG=a�t&�c����G>r�
�����t��h��az��՚5����ި��)M�2]G�K(����5Vvd�ē�6�Y�Ď�ͼ�8�.vDY~��Ks�-2`I����Vlv*�go�Ҳ-��F�d�f�?{g@П���Z���u���?>޷�U�p�~�ցd�������$ f�Ⱥ�.fx�] x�X�N�>��s��Қ�w����g+�N�����>�����ܷ��}�4�t�
ee���)��L��vY;��äͲ�j���z0�8z��m�G^�7����Y�Wp�o�m'�Y3�2�4t�p�o9p��έ��)���90�r��R��J��'qƘm;4par�`��U�i8`�q')xpƬ!��v,��h:�~�q�мf̘�g�'E ��T*���>���~���М�7���&jŲM�r�z�[T���� l��[+m�i��;�ENQ�ض�	�d���,������5��<�cVX0 �M�K���1V�����+v������x�����{P���3���{�t���9�+6������;�>0��uv��l�*=�p��][�>��;f_�K.9C������}���i��7�;�ao�r��a�M*�����r)v\�v�j�oV���@إO�`��ybY1�#�1��<��.��0��8̔k�)1�ơ7op3���ǎ�qՂ�bω�0�R�+J4�B����`� \Xv�� `zY@�܎�t�[&���2O"��]����G���Y.��eĪ��y����Թ�C��{���(� ������g��eK7�]��T�֮j��n��}L�� �΀�ϵ�����x��) ��o�a����l�f��2�HM��g'�#C�K=��\|����"�������s�q�������̹�;���|cv�/e�kNh�������ڦ��U�5{�.��Lm޴I7}�.=��f�s�n��^�w�2#���Xަ�Ɣ�lWQ�9�CD��x��ؔ��31�`�6�`���'59���qm�o\ɐ��T���
ګ�}
��^wۑ�����jI�".������	�1w��G�XK@�Ѩ�P���Ll�r�=���6Qx��tU��Fx�/����ĽB���#x��Ȅ�ӧ�4:��:+��f�}���K1�@}�ԡ��ŋ�k��7����0*(�p�c.TQ�];�\n����M{y����P.��?Nրh`�
��7����6���r]7!vJ�m[C�.�3���.fb��eg�����
��;s,�a�1��@�1���،gv��0�=y�@�����X�Ǿ�@=�4|XBw�}��N=G۶l�'?��?O�B���ןt�&w�����.���T�ϟ�9��V�g�uV�%|��I:�EH�&���*~�6]��
���́6IX������+�x�o
��p��/��?�V:�P̉>�m!:"W�Vsk��1N�&�4������fR#DK.'.�j� ��kw`���s���XQH�#�"�ŕ��������xІ	V+�\���wݬ\n�.�r����^���j��k�+`nQ�<u��7^rPB������`��c>�D�����˯���8^�}�c}_~�
������]:ۋmZ��$��企�lo�lw���-�8raW�tO��33���	{��}q�.A8Y��K5�#*�t�m�t��4m��x<�̏�K���ϫXn�M�Cc�zk��L$ECM�|��ɺc��6�c����o㋽�\�H!| 4c�ӟ�t�W����^�r.�?ĥ�L?��+Lp
�φ(��'��g3o9�5M"&���y���e/�W
'����\S��.��l�1�Mԉo����B3)�1 �d�1��7��v!t��Ht�����������,x��~z��E(������}:ċ���{lی ��u�?����z���*��V�\֦E]p����;kXKk��+u�Q�ao!}�^Lxg`3[�#l�I��[���(�3��Td{q��7��F9:���!�A�n��b�pVK����_A8fJ���f�x��&�3>�M��?�Y�'����p�utDM�V.����/��-�[o�����U[K�:�KZ�l����s:f�)�d����^B�j!�Q�^g#�	�NoBxΛ7/�ѯ��}�帆﮾��0���6[G�x�ސ-I=בI�8Nn�w?����0�܀2��duȜ���w�sO�{ｃ[�}��|��Mk���r`#J���:n�&O�4�5��z�kO\:n��@3]w�F���R�� D��sx	`
�E{}�������*0�_��^�Č���5aK�n�uޑl�7(ky5d����!�Ӷ�5�6�Ce��/m��_�B�AU�Bմ��M�RG�=��~��� ���۫ /�̈��_�r1+f���Px1�s�u.C�����D�_��#ݛ��}![O|�W�Ǡ:��&3Ƹύ��Y2߹nn�t�K��I�q����jǽ����@���Ym��HT�l�-\���;�jx[Vw�y�&O~��U|ERcS�:��Z���9٘!�t&2n�[��l9JYƊͅ�0E�w�y�}B*,w�����׾D�P����c�g�F���1�l�u}�wl� �7���T~��D��H$�Ycp���Gm^;����6��ՊԚn�ȑ#t����[�<\���9mܸ9h :e��
B�|BM��}���q�&�Ɖ��6��\�i�L.l������~��9T���k=>����=��Y+(��Ѷ��LKɜ2e5-_�]���W�6��%K�ӧ\�qc�V:�Pg�$lP�g'!j�����p��
�ūgG1m{���I��]��w���cQ����������TzE�?�0fz1 ǡ��x��α�|g��ګ%?�J!Ί����
�^��db�;�=sĪ%z싏*�ա�mM�|��:��w(�%�?���(�fK�����$�4U�i��0G�2��~�0'xS Lv0YL 8�#�3\��?��`^��	�ZVvA�ۤy�vx��5ϣĀ�R��3�J}u�w[�GoY7�9���D�sò���t����굫�Ң%!D�F0�A9f�Ih1j`�y�駃��n�Pb���g�}v�� S�?�q_	ź)�\��2�X    IDAT@9m&Y`;4z�ZT�ܭ~�_�e��P��L�j%�Jy�֯�R2դr��Z���UM�2K���t2[<�w�;[�ƀ�h�]��}����U�d�oX���۹����-�����@pꩦ�o�ݫ�	�fY��������
�����n���1��Nc6(�~|3�o�
����_Z�HO>�
�|�H8��U�ښU�w���g�E��S4z��T����O��a�k�U��W��v>[a�'<�|�M�b �܀�9+�&H��"Q��b�\l�3�����e��C&|Q����:��>��~ �<\�����}���!j�L�=�#�V�P����r��k+`�%ځAb�o6��/ɻ1���л��J`u�%xY�J�_=N0�jQ�D i@��E�=�b�SJ��[TcC��96m	EH�	v��	�w����
���O���`��'
�=�<���v�>|G�aL^A��v�mF�Ն�ӫ�����A�w��]k��� ��x0���!�mG�kT�p�!ż��n��l���۱+Ξ�#��Z������խ�tF5̉Y�6�R�*j�*V:^�)�*I�%=�L@���U�Ʌ�K��o��P��F�]�>�7laFr��3�-k0�)l��X��vk��W1��躐�ìA(�O>
C�,V�U@��s�νip7�����#7���R�>&�9��чh֬+�S����j����`�A�F4ڱu| �l�6��BC�N��`8��s�	ڎplϘ%0e0�|� �y���A�~~�ew��\T������B��v%��'WS&�Q!׬tf��h��.�eM�
c��1s��s�*��Tcd�l{��cgVe��5��U1��펾��ڸ7���L�;���<ۀ3_��ݫ}��n,�X�Y9%66),��8����O ���Ήw�v��/b������x���{��0s+V걅_R��G�DM��6e3 k��ʨ��j�����<\�dJ�f���3&j�@n.gi�1��v�m_(|�s,��{�E�k E�E&&0�|�6��{G>�]��^��^�3��Z����o}K�j}�@8�zjޜ�T&Nx��� al�8�ƿy����*=����_P��ҫ��p�1`�DZ�P�`ԟ5X8;/��'��h;�'�k��&����%�k�n��>�9�X��oK�͋E�|x�9�C0�Z5�bn�~��h˖5��ra��d�I�|��.ݢ$�Oq�%s�97}�e7�(��^		u����&>>��g�"J;]��Yml汼͢ݦxij��g]�j�h�nWv���y��f�՞cZ��#O Z��Vef��x�j���6  Kq���{��7�
Kwf�**fz�{�$o-_�Z_����uu*�(���M5�;aӃb1����\�g5�ua���sy0}_Q�|�P�����sa�l.K�m��"?�l�!�L���k�{0�T�՜�1�����J��^�rh��v�S�$��ٱZͤ�_���9��[�='��|�	�8�m�2e�~�_?Һ���UQ��8�H��e;q"6	`�A���Ʉ��B������ H�~�,� �ܹs������߅R�/����c�?���h��$s:`L��s�C!�l��_آ�n{@[6W��XJUKV4m��z��`JKb	�e��}���~�~�V`\g���o�|�X=�|����	���N�ݱս��1�}�l+�x%�@�(��\��8��e��M6Sp�:�*���}ضH�0s[��"���2�\}϶a�Ǹ�� c�s�&�zD�����]�)�]�A=���/{g�wU���]g�Lv�UYٷV�E4 	���
QDY�E����Z�B
T�.�V�\�hA\ؗ���$$�}���~�?�p�w&�dk�:וk2��_�y�s��~���tw���m�矡Y'q�`?�g��Ʃ����^R=[��|~�����L2��eW9��,ކ�x#&]�5!��"���� ��c����
pSmyĆ�棵LL���B���;{��%#S�j��$��h4���}W\�ы�����;c�m�۬Yvg{��P�lX���	'�E<|�֭_�j�2��V�a�µ_�:K�P@��\�a���p Z,�����ٳ����a�qx�OX8B(�]���ج��~��5( RR����T�s��պ�y�K��~����������k�<�0 <C�75����k̪���1b3d����1���f�1���m�ɏ���A؆(��l�l�F�G�4p,��F&8%Ly��d� Ą�p�Q�b`Hb�f��6��*� |��q�et���@��������>�a�8��%r�a{fɳ���w�&�e����B��z���n囊�h�:�2Z��/�`�U���Ԩ'��S��L�a�q_�Q�>餓��#E��z�	c+�Py;��
�L��0(�
��, ���W�}�,a�p��kO`��+W=��Q#&|͂�;찱;ވ>۬}a��Ca���3�x�	����*0a�#PBvj�v�Q"��'��}��G��k_��`�m������ �2�����;/�7HUÅ3���s/ ���q�W(���{nծ����9G�e\����^X%�z�T)OR����蜹��mӶ�1��%~5]�6�R3��و��04oAgl1�\��צB�N(�3��C�(��PF���CHG2�i���|�.�B� @�>3�a�� `�=6�iO�@��a#������
8����=ٸ�~���"��T^0�]s-[Ӳ��ۿ�j�&�gt��wi�i'h\���ݫ�>�L?��ot�NҤ�;)6����2�����Q~ I��:�������pe
HiE�+Ű���½������� n�̡d�_�	��˹�������g�;��5�S��V�\��]{��c^�rʺ�'�ˇQ;�z��춗�<�=��
����z�,�a�q-����\�b(
�b/`�-���=��&fl��k�b�$V�1(9+�>�Ɩ9v�`u�����2����e�]�re��~���я�7��=ۥYo;G��dU9�)+�9s� ᰅ.)쾙y�[���� oW�3kq��<q7�.�38b*.�v�7��"
rT<�_���/ڋ~9�;�}f���"�O� ?���7���'��nﲱ��6h�͌��f��\����������s��v@V\����3?��Q}��E�'�/�×�Ws�Y�J�~���u�u�V&;U�/�V�L�_Ŧ�����BzA�L�~D[b���7�����v�ϥ���'�0ǹ����d��0@�X�zꩃ�`�Ƚ�,��(e26�F2*�q�\�*����Ύ�Ps���c
�u��v��q��ÓڟE��v�駩yBQ���*��I#Q���q1�:��RlmF �hX�?��?�O~�q��!�j!t�q��^��,qA��dל'��]c�� �(uU�L^=�}��k��C?��{�����N;３��J��K��UTU�h� �ʑA�<���A�ƌ2�N���%�ڟX��1�C(7�I�7�.^C`�1a�1ۦM}?�^�H��}mⰾ��Ô�P�d��z�Ā�
�����L@L���sx©\�� .�|�O8�g�p|?���>�)�Pr�ʗ�铱yy
��%O�w���f�����|�9�M�бZ��S��7�S;l��.����^*3�5j*���U�JJ_���46��;��oX�SА�7}���?���&������:+�^3ރu���$���+�c<���8$��n��,�J&i��\������c�S֬^�V�=&�f�u��o����/�Z�R))������U`O,'Dc�}4;��VpPRL��ߞ��f)o~�C�0�0
������0�T؋�,:8���Á0���;�OިG��c�Ol�[.�|bX��~�zzra�rEQ.�}�W.07�Gl��ְ�?�{��� ��xO>@ȏ�c�Jf��b ���+ء�g]yW!F�%9}�=%��c��+K���Ϝ�����9�.p�qh&[�z�ސ�5�VZ�jc�}�Ke� 4���Oq1����\!���I�FhP���I�� ��h�%������jG\~�_�z�ŗ\��=��&N�S�_y�v�c/��P}��W�a`ja{3?1[��#�<*(y��ؿ�����%�I���<�`�@'g͚�@>L5�#��F�^��1�`A.���ųY�C��|�� �7�����pјo�s�k�.����������O�v�q��o�;�����Y/��X���
:�%Y�d+ ���"On�<���qز�\C���?�?Z�h� ��� R ���9w�DҮd�)��:_O?���͘��}��`=�||���=O��#� �`�3��HU�6w��O���X���8����钂C,`��Y�</�{�_�Ťe����=�ዑ�a�3#�k���LPқ�2��.3.o}u{��i<D��Bs���t�<�m֍�:���c�f�2 /����\��szn�
ݵx�*}���.]v�;����^����O�G�L��T]����w��P%��l4 /���,r�&�0?�H�͐7օ c�kƌ
��#���w�uW p��6b0W��3�fԮg3`�o"���cH �9������Y�p�c�S:�_���uDH�md�� 4���o9JG��Z�t�{� �X)�rc%�o[d�8�@���.=�oߏ�8��E9��(��Ua�U�e|�M7�ϓ�yIa��03a�>�eg�������J=����y����?+���V�\��k�aa�Nv1��9M�����#�ir�O�Y�Ȍ	c#135h�l֬8��oJq8�L��w���7��>���9�q7w�~t� l&N�!��Y�S�b`��@a����j�fo����6��9�#m�� �������)�I�ce��ιD/�[:C1᜖/[�;�r���^��Vt��gjC!��������SWW���˴�A�+�e��9� ��I55)���E��ǃ�K�/�����
� w�_���<x`�?���y�I���FF�����t��4�����>#���;���f�s�7^0s�̱ˎ &�Æ�wf6�=��OkK��e:٫v�NG�F��k���\��6���n����R�!�3tP�+�TK;��#�p���*��=��u�-����}H�'O8Y L&N�m�?��{�u�&��Q��)T�7i�ҪN�s��;�Tm��N[&;b��M�[�|%����o:Oxs'���u#�Y��8�O#���I�m�q�5f�CńcY86�g�0��O��z9�K��m����7֛8�����/�F�����\됆C^���q���G�����M`םv1 0p���} ��h�.��p�ւ��+V�+�~I�r���}��Ӗ�<VM�eut�����Z��_S��	S�U���,�ǩQφR�6.��4U��m��c�]j|�f��/�8x�dE�u {�Ћ�>{�t4v����"xl~�z�9k�!���b�.19��d�{��7�o�AxʚUw��&�-���}5��4k}�:��N:�-o���3��E�⣋�披EpD�)=Gp�!:��3�;wnȂ`Cq��|�ɧ�ӟ�tp�H�p+�I�r��0�es� ҡwh�6���ӻ\'e��W�ӏw��9�T&�٬Z&	\͙�A�{)�gQ�:���ູ�	�q{af�N���� h ��w�@g]2�3�t@����e6i����~�C#�g86S�-��Ôx�/~����Mq�3o��
d��q,�m�;��o0C~�g��]j>�����=\u���𙋔6%,�nݚQ�0�E�s�����+�>G�N;^��z����Fmmؘ��5%e���/��T��X�J99�֍�a�.eI���O|�t	9��w�������B����c����c�l��Ϙ�a���Y!�l쩠���F����r����d�)f���RO��CY6�N����k�����;�J��7T �Ӗ����i�v־�N�0��(尢�` �Ap�k����i#f�qY�$��u�[Hb�(6��=�"V���cΓ[�0O�֮c�KY�|M���6�j��N}��VwWC���ҬZ��Sg�����G<����H`�%��t��"�}��w!%��x;퉶��f��JG�'�}L,�cc���ص
,�F`K�{O�7^ȏ�]�!@ ���3���6
���33�o�_g
��.�E�c��$F{ i�0�z�F�s�{�k���X����>o
��b[��1̗ԁ�A�ٌ��|^���e�F(�_�k��x���d�IH!,�LP��I���V4i�����!��d���,+bۤ��xi3&�Z04ȋ�g���%F�c��� �C=4Md�z!�qhgz!_�1��p�����0�_,X�1a�&�_�#̄a� av�UJUm�������w���	a�Pv��k7�OO���"[�j�&�$��L���7�'��d��n��"A�ܩ_�Ǐ���uji&e�'1�f=����8�jU���ե9'�����;}�e�-�?���:-9"_� �d��;2f�G�v㝞�1���=:D�p�ͨ�<Zy�G&6��
&,��o�Hy,#/�!?��b��1Nڊ�a��nב���gB�v�����6�@�#��i�`����y�Á�#O=�yµZ��Ld} '�Kjd8ȳI��6���4~�P��y����F]��a2$�!�D(�Fǲ t٬;G�;r�%B�����i�����'�`E~ ��s������l.�8��
�x��ⅹL&�ʂ��p���f�	s�'�lM`�J�w��p�*I�C���� jf΄$��F�q��V��8�Y�cA{Ų�U�B%�Z�[��U.7)�oQ��S��B�Rk�z�f̜�l8i#Y���{F;����GNL�H��zB���8��8�h�06ncNXw�'���X�F�n�J�C��M`�Lf�D�5XY�&=�3ș�%�IL�Ek@� I��A�n{�6�a�� Mϓ��� �/`��C�m�	���%?�qzz��}�=�\ߡI��U+�(ñaY�T!\פ\�5��q:;�7̽z���0���f�p=��|@�= (�A&��K"��9|�3����f!#dF!3���⸱�o&< ��]s�5�9��~�m��#�c��<�1��Yi�K�"����PP*�:l�	%wƅ]���}V����|��SO����5���W_O.�P�\��+e劍~�s�Nꡪ�T8�O���0<n(#��$wZ��*��s=Gۯx>�	0������*�0ڶ�~����	�X����X��۸=��i�=�x���quH���L(�{7 Y8��3&�K0�a�a���c�����f@x�[Lyi~fٳ�����b�Z��U��J���y�T�*[��n;k���z�31�$�!��/��!/���CQ&�$���ymo	9y+�=a�4��������2r�VlD���=�=�rc��o��׭Y�^�=b8&#LO>[y�+�1���H�z>� ̖�.���0���v���K�A>V�F��J�[?�����g4���<M�d��_�bq��J5�
 <�Wف�ԯv���)!gLw�,�r�b��X����)�Ϫ?���c`L��~k�wS@�w,ް��q���F/�ŋ>gB��8��	n�Π����]_<�u�>�B&�P�<�������;�._�ܨ%�̼v�)6Ȏb�˟5�{zU����o���&�+����/���=�~���q� ��,�}��I=��2����EM�1����X.C��-�{�<��X/N�����j��L���P�1�k�\.��k���1e��׼����7��0[Io�$4 ���%3;���@���Yn<��3:O,Ѐ�������ꓢ�#�F���zC%��S�}D-���>E�>ݡ/����    IDATJ��y�W����5�a�����CHt�3����"p�PL��6�CyE[
�ai�	ב�t�K�c�����0D��`��&k�svv�x	��p��U�gx��Yxy>���x�;�`�}�'��X���W�?��7� ��8cǼ ������M��,��dɬs(���ҥ���۔���ڒ��Kޥc��3�l��H��/��Tn����q��T3�e[�� �/�^aQ�� ��`�l��cꐏA��3 �X;]��}޸C�A�`���M8r�ܿ]s�5�" �V�=�U��1�d�cR�Ó�V4IKv���`�.XZ�ce@x�u�Q@��;Pp��k; �"Ύx��������zVi��NRKKU}�u�x�����is/ToO�JՂ
MI���S�j���+��&�{^�1a�U��� @�:f]6�1��R����s�����>�$�[9V`<��3@ ��������	O ��kv�N��]XK������1R�.���j�T���g"//�J 0l��Y�">̵,���!���{��_B�rZ��y}�/*��Qss����<�:�8�8�F�e'��?��ϭS_9���I��,+�mW���z%�}�=x�v���]�*\����c��A<�D^�C�\���z/�ǀ�^�0y���^�ך<nc���l���]t�n۽����K ��J��Ϻ
���՗\[O�TS�x0cv�'pz���y��E̼�!\����f��ٹ'hF�u��O�-�f��:􈽴��U���:����vMF�ZS�X�f�</l��e9$���M��1 �S��
��-��0>��/v���r�7�o1�<����I����c�����h����z���AO`������ ���y&>�矋T1o � �k?��={y���e ��s aV���qX�g��1>���%�>�&�՞�e�� �r�*�~ۗT��W{[Y��;4��7�ؔQ��^������|Z�F��^��]�ϵ�\��X����~6����#[ד�m��蓳Bb05��`�޲u���!�� Ӎc��t��+
�ۮZyW{�/0a�3I�0��3�cf��'��	Sw�k<��'���v���oTQ3x�%�8C}]r�{��������U�/=' �SOn�;Ϟ���R.	�d�Y�}���"Ȏ0�e<6d�ԯK+��(��`4���c,��cθ�~@hF2�c7�^�3�T[2q��1��粓
0!�ҋ��V��d�� J��H����� ����Ʊy�c����r��llr�E���DV�1X��X�c�5^$%"a��8&�iC�ӳO-ӽwߩr�[���v�	�J�O���[�U������aG�H�}��vI!�I_8���k,��	Wz�ƞw�k���C#q8��3����r1�dan0�0L�l�\O�v����t�A��wbS f&�8��<ǩ&���	��H.���C�/�ȫћ��_��~��������w߽�rEI'�:G}�mR�5T|���'���f��ˊ��qrR�; ;����d'�V�t��bH�hDf�V��P 3b�,�|�&쉵5r�{	y���[�E�����D.�8}�3>�6���͡��A/$�� /y� �]rX4��&%�6�� p�(`� !lݛ�_5�L{�U2�rZ�r����ڰq�&���kߧSN>>��-�����2�膅�=����4��3�'dP4B�D� �Y�Fr,�'��=`���A�u ��M��rp�����.}磌�:oLO�skW��^�ga.�?c&�UR;!m=���غѱ8�.fR�	��|}�J������
<��0�E�;�Zx�U��#�W넒�|�Bx��z��:������)�[��S�N'�r�^7� ֆ2��D�)��L�?�{~6l�9�W�c���C�n�l ��Ӌ�2 |f#�1�.���a��O��X����������C����0;�`�;��da��o&?!<@�����=���;@����p�����l$!E�8mlH}dǨrz���oܫ��U�<��˯�K�4�Xm���/�F��2���?�j��?a�J�^U�%������4��Ĺ�c�A�n�����>�(�XZw�=��c]6��׫����1a�-OzaL�s/G�Y���Asw ��y�o
��~9��-��CV�pލ��x#?�e`]/�s]�n��Z=��O�������ߠ=��K��a��>����ʩ��4��P;��SN���,Ւ����WyQw��^�0X��D+}<�caP�X]���+q4C�#f��9O,_?�e���;E&L���a��S����v<�� U��,�x�Ӽ!�qd�7��4%�IZ&�)��8�J�:�@jZ�g+&!6O�>�\�l����E��|^�ƕt��h֬7���G7��	O���>���w����\PWOg�?C�B!�$���nCb�6q�o8=2�ݔ��a3/��ld��%��t��\�y�r��.\���1-e9����x��r�aÁ0�����]��c�A72�'��C����5�\�x��B���3�v�i/�	�n!1�Z���?z�j�U:�o�g��V�g�u�POOa �{>����C����B��"3�E!t<����d�Z������G��ً�+�|�p����Y�B�	�`FmX,����E���/�]�>��t�� ��<p��ɒ��]�B�qo�u���v�����'ǁ�qg5��|aT��w���s�m��oPss����b�|��d������?ޭ��Ї/�V�f�l�(4)�M�- L�i�6<V��i�I@�8{����vl�z�U̃o/\��}cz�F8����{u:V�'LL�ě5L�T3b3��:0T�'�n�y��<���B�e�|O��pD:&��S��>��oi��:�35uj��{���ɲ�<=b�N"��#V�'�3�z&��11f��&�P�nk@m$�{Dą�o'��<��f��'N.[���]b�.a��a����~r�d�m3�r��a@��7�:�d���=�F�v��]�)� 2� �yƄ#	��|��9D��C
��.yN��M�z��Œ���/u�)Ǉm���=��J=��J��4�����96rp"M���|���a�� �##�����66����8��a;�wa*/�zm���#�s�ܷ������9�~�u���!#�0����
��������B���=1���-O��@`B���cP6X�r�7����8;�q�
ɰR�Q�nפ�vjҋ�*��W[�6z���:�����ʐm��:��5t��yz��
��$=-)$���y,�x��A�1 !�ȴ���X��.��G����?ވ3�V۸C�gs�֦&?�u.�=�V�3�+�b�Q�7Ġ�^F�x����D_��ec
�dl���8LF�_�%|P.�n�;�q�pQ߂����K��2��@�*��زH�khժ����I�r�&L(꣗��S�E�:E�
ji��Ξ��[�J�FA�-����W1?Q�|�*��"���\wi|���3��u�{\�1��I���PQ���qaH�C$�W= �ߢ��A�����M��|��g��eԎ8� ��q5�#��~Ǡp�Ր^cpuz���t����W�bBL�=�0�p�����3�(ꌠ��Y�����7[4O9�A���a�TQ&ӭ^xF�dU�_�b�-Z�lI7��yuvV���T�t�����9� e-I�ګ���|c6ʢ'qa&w� ��cm� 	�2i0Ƹ�^�J�Gb�ǵ%�&�W���'�}<�@X�� �	@;Ǖ~`��k���o�8�.�@�g��u���ʞ!l���dC�>�o��!D|V��Yo�c#~�K!�Ax��%�p������>�zӛ�T�ҝę�ֲͪjm��b�8���a3T���ib�I�=�$�h��6'�5�c0�G6)��qp(Ƭ�G�a����wv�;��s�yޥ�N~q�ɍ��=�]a�!�J�,RԪ��fL����>v�hs\T3$ǁ�������Xx
�s=�q�|��'�|������S��T�{����˘�(G����xw��(mz2�uU+�����]}}T���">�RC�R�::9i�|�lO؜2w��|�5a��$�$[�_�?��qYD����4��e�͌f4rQ���opӃKY�
e#`#k�7�`$wכ,�61��G�"�!�`١�a!l��6sX;��l�� SH��������~y����Z:r���;�YI^�p���"}�Q6TQ[�b�����HU�!7�6�O�m_ԥF&�RoQ�ﰫf��&L����B�����dיK�z��c0b����7��x�	�S�X�d��xa�s�%�����H�Er��k��g�End��0�T@�Z`��{3coj����L&�\8�Lxƅ�m�v����(`^�6�s�zM�BU3^��������>!� �ԧ)�H�Bh6�Bz�:��@3�u��t>��yw�q��������PV~��o�&�0�c�9F���g^v�	�cZi�|��!$�У�>�Ro�����^M?I=]R�i�*UJ5�l_X��{�ٚ6m����X쓣�^�?6`���DQ`�;p���w��h�³�*�(�C"f��-�4@��|4��^ރ�xLlBo,|yK7zM��v`��d�9�� ��3���f `��9 �x<��x����`D�`ڃ�nX<�ט�,}��{:2�#�>�;ݭJ_�*�t��U����q�p|Q.7A�}d*�IS&�yCK�=�s�0�I�tE4�O��	�����a̚����� s��� �k��
+�'�`�]�ݞ��u��`$�4���K8 f,h+����˵�^{ј���,j/��p��b�®{����6�Ӳe+B���h�M�K�@�J"4�]g��5 ľ��m�Q�N8!��}�����gs��fፓ5p�-#�;��#f��3U�to���K����~�Ҫի7j¤mU�g9S$Z@x��P|>O�N�}u�178%(�A���j}�������|� �DcB�v4�Ǡ�c��Z��L�/nͻ�r��8%履�#�it]d���iz�d���M�H��C�`��9o� 0I�7��p����w�6��� �P>r�^.�X'�����%����kɲ't��U�mRS��\�W�ҋ��-�*�m����@esM��	ƫ^�"bF�}�P:Y�\�+��8:��@��tµ��r�[�s�}�7�ac���H,3��ZF�6�`��]�1K�����1�e�Y@��c��_�hۜ"��<N�jV��m:a�����{��?@ؕ��xfE^0�$!4�±���㸕'2�b���s���(�u�]����x�_+������ٸofo1��چ�*�6�_�s�:7vJ�����sEe�mz��U��[U�$i4� <}/��Ձ*jM��R&l�4�dl��3�2X�<�1ak@o�{̬�Έ�7���x�I@0���ۣn�;�>�X0�	�9�H��l	t�z�|a����:˖���?�i Y� �ș�p-2�~�=�;w�0�F�VM�
��f��UH/��?����5�vJ�JI;�8A-�R&�d0��8q;�|���m�}T�'������{�9R[ɰ���y1�~;���81���w������'�3�� ֐5� ����*{��g�l�����³����p�C��[�^��r�o.X��c�SV�^4%S �i��9c�~�5�Z�f��z�i��&�B�*!�3�!�V\��N��� �^���{Ă�"�&9K�$.��<�����o���ͼl�`�����o�)_�R6ӣ	��U-w�����{d�.��@�	��4��>��|~@yY�|��YO�f �ǘ$� ?('���΍�lDc��g��@G�0,���Ys��Ѿ{S���KX��3�&��	�sl֠�.X3���C��i���y �s\�g��\W��0b��;�U��)�#1��K��60�'�zT_���j��j*J�;O�f�\�B�v���ꮄ�����h��ev�����)��2����A��L��+d�gȒ�:�$ ���y>��@,���:gW�5��N��^̴�y>�s �{�'`��Q�V�����r�!��D�6��pso�A�����+�SN����_��~ul������r��s�(��M����(X���ٚ̝o�2���!��8���dG���e�	i_Ҷn)�N�nۢ���ɒ;ث���z��:y�{��פ��j �,���|.�W���dDff+�9ed�����-��a�5�y���5�d,y?���y�=*��h�vS�g�qYЁ�B�K��d3��j��/בֆ�9����@�(I��x�f�qxs0�����s�s�E>/p&��49�Zn��g2";��/Q�>M�ׂ�.Ҽ�OT��Rؚ[����auu���P�S����d�l O�s�v�X!/�
#�#p��=a�#�u�r�l����N
�x3�מxD��.��&����7^�䏐���Z�V���},�xLA��)/>������B1�r��ݷ�U�z�;�b�Z=���b�1~i1��Sh��`k'?v]qP*,44�ů��\���Ș �����Ზ��<I�܊��X� n�У�~����L�)sߢq���j�ji���U�o��j ab�a��K��pD±��@�UL>����B��N���l<]d�c�:���3y�R��}���� ���@!䙢��a������:�݇��aa��88�y.a<FdͶh{0~;B��q ����Hy�=���l���m>�b����/�V����u}貳5{����e���o~L<�f�8R�l���
;�Z!�̚
�E�O��zǜ�l,[���!�����!��v�w�y��w�yg��E1�1�d�<`������_��R�����{'��"]]�֢j�|���^���1�k�/������NJ=h�:�y���%O�t�#�0�!�Kh�]4&�Y�Wym� �\-r��c�y����F� /l��o��E��{b�P�L8��V�z�_=�kt�՗��g�N>�X]����5�G���y���E5��x0�/��9]Ӧ�|XGxɅ{��0�J�Γ�c��;��Ŵ�ٶdru�W��Qy�x�:���nh/`mjG�h�e�r�����β��i`�,�՘�S�(�ü��0�a8.i�-�0a�8���c���N:d�35�����d���Z|םa����U}�w�3���?y@��?j���.�kM�v��բ��%�^V6Ǯ��td������aLa���1�<�G�Kb�,ԓ����O�!ț�8)�5�9��)������Ż��l/�﹖�ID t��3ٺ_��j�|��kn������o���ֈ�5&�Z�hJ�q ��t�̃C8��?�ZK�?'��BH�0�
���;n��P����.��� ��[ɉ��x�A�l�@ ���g�pPZ��������p/��@���(p`x����_.�u�]���zXS��붯��^��nz��:�B�F�\K�u��9�����d�k>ʓ5�I`��} ���zP���Xm̈�DF{-�i��88�?�b<��{<�}�A�߱[�^�L�O�����[��v/��3& O�u�sp~�Cc|�gH�&�5`���x����yq=�0��L�|���-c/�� ��X�hb����V��oUϋ�0���^�N�|ʛ��]�5�������4i����G�����U.OvUF�ZU�BN�P'Y셩k�I����J������Z�#;X��?��p�����xA��~ثpx�ޅ�:��K���݌	�;2��}q���E��W]=L����~h�I�W�9��H�VUԎ8�0�t�,���/�n�ZUJ֓�5X,2|2�����ut
A9�������v�m�s^q�3 �-oyK h,��,>���0g���_�u��9vcE�qa�sl���S��c}�n��:=��o5~RC7�C:��Ѿ�q5    IDAT�uݚ5���4����Z�"'���	�MQshd(F2�Lw����l(��y�E]|��~;��+06��\��㉀m�B��G�V�5}��I�3�aY��x?� 8��6Z�M�v�g���.f�<P%��� ���qȇ��0ۀ�� �2�ŋ�[�+᧟Z��~�N�z7h�Ć.��,�tқ�am�.��=���~�}��_��4S��b}	0��/���<�f]���g��n�A.0�P��s�f, Ɛ1Ǔ�]���3�y��X��;�;9���	��������6!W�AX�b��֔����]~��z��m[�#֯�����P�Y�����ЬYoӯ��־�F}=����D��d�B�,OPB,�58l����ɂa��
�����{  ��Ib��(��t=a�3a/,�)�ro�nXx�~�˟��Cv�?|�Z�v�]�?,�9�H��Y5���
�e�� z@���F�1�RR�g��P�?i��f��<�q���s�ꭝd�N߁�X >c��ǘ�۬�qf���f&���K_gC��5{"�`e=�6
�k�x>���c��aWN��"`0��.�,�9�3�7�^�Mf��K�¥��\sD���"+��a�n��~���+��[յ�M����׼S�g�Ύ�n�����>���t�?�LW��)�Y�(�YQ!�{��Oh�e�¬R����w�;�l�r�3�����_���s`��#L�x6^��+��m����Q�QJ��"�E8��R�T-�͎=����ի�l+��R�QML�p��5K��G~7��!�����e�QB6g�BƲ $���_���+�8��ěY���e�vBA�4��+�NU�~��>�7k�LC}]���+�ѹLg��D��]�B�ӧ�\�s���[WW#ۢz-�l�%���
l	0��9�h���Ō��,�-�}a���e�¦fh�@����� l���^�ݢٟ�x8o�+��8�c�h����6Hq�G���{ ���g�5.$c��
=��X@c����3/�CΗ'���x�KtP�}{�<q���sk@���+���;Gtj|{EW]��r��[�������S;3�����}�6>I'$5�yT#S*I5$!T�_W:s�~�h3��
���"}�c҇�c�`��@5A�x+`?f�� /d�����H[�$Ƙ��?���z��"u�\u��fG����z�0����^����[&6���ab���7����<�(n�­ fC$.�LV%�w�:�zK"ʉb��0���IlwvĐ1�lM��F=��/��n�5c�.j���J���/��Yg\���&�5esy͞}�f�<0� �誨�Y�A��O6O���dw�w������k6N�b@J�S��H����i��h(�m�=�Ѽ�F����1� ��?��\�F�UG:/0D� �\m���p���w�AR���zb� p8A��G�M���#��Kw��ԳO讯.��\����L�r���e��k�~=��M�fg5�L
�*��Z��ve�lEO@�m��$-;"��q���n��"�	P�Ff�;l� 6�,R�LҐ��W��8��s#§n߃AMy8����1jGd��o\;�y�1qՊœ���j�Զ�zӛ�ӌ�����Jk_X�r9�c9E�Av�項���a��A�X*�j���b���ISC���$@���Q:3l�-�}��/+xb����j���V�.�L����׺��7��?��9���֯���mV��JnA�O>}�	'y�c�3u&���m�c �Cf�q��,4^�Ќ�6�k�׋v�o`6 ���e8��6�n_ړ�e:�$n}R?$�?cc7b��È!+Μ ~K|���`x '!�+@���6{�{��\�Y�?��p�b�̛0 �}�7�K!=��?[��.}*d'�<R̕t�U��ig�Z���T&�$�V�Xޡ	wUOO]�zN
e��jToY�<��x�7�����S"�����~7l%����L�!�a� T���K�"o��%�>1n�'�
,�X@�@��6n����������������ï������J=���1�L��M�Wo|�B��}B��	%g`mM��v\ǹx(�! ����ʧ+b�Z�LB
�\rIP0@څQ�Id��0�aet\��*�'z:~����R�Ӓ%���)�L��j�S���YU�7�����%G�$ LLx?e2ĞQ�х#b�f�]f�˓� ��.��l3�� �H��u�&�A������4 z�Gz�pߧ�f�N�73��P᝭iG����{b�3��x���a~3����N����u;���E&�8�Cx�� ��P�Dr��)����D���۾"��j�Kg�~��p�~�zT�R��MM�SU-OЄ	����������JT-l
���-s٘apDGX�!�@H��0^��g�&j�xӘ� ;��;����P�u#֙t+ި搩A���	<�ZO�����|.��k\;� �M��řkon)fX�ʔ� �qo=F�gLӒg��s�%q&�h,�`�B�3������2�ʈp�^\CHdF�
z��w�+��Au5,��7�blN%��`N��$���l�G~��֬^���^57eB"�fM���mR8����O �IQ��ד�)UN�3c
pܯ��-����l�l�=q�y�-\1�؜��k�kE����������h͜<C��t��c������
g1�m���/\�3`d>8������8v�wZVl�^���m?�c�2���z5iG���u\U�q���	z�Q'��}�s�������|�/�-�jo���W�#�X|���h����îC�+��G?�YT��a0���q��
u���i!��~�7 �aT���F.��Ƃ�_&<y��w6uo<&�Ԅ�i��l��O�*��]�b�։N؂��C[r�e,
�c(B'��vĖ�g��F ��=B5�5k��G���␄]A��1c�|*K��/�鬫Q�(�k���Y�WooWOR�2�d
�,��Ve0����&��هc��,��@y��o�'^��A(aČΟ{1y�/�,;������K �1�JV L�P����F `�O?�ϙ;��Pf�\k���/f[3�	��e�t�w�^Ω�H!��IA��6�z-��	���λ*_�T�q!Lx/��7��$Ԓ,&����|N��?��C���� C�ϟ���7�8���>��]���ο�R&cY����Nj ��󦒚��s�V�5�-_4���V,n���/d3l[v=�Z������POx��v�c>N���q,��1+�)����)1+����b���w�3�����Rc*y��6�%`pI�q�%��%1SE0��>�J?uA����
;x
M�/T	���Y��e4w�;4m�tr�Qݛ�~c�d�n]ş��nc���$�g�y"�8�~����������@<;�=5��F �����t��t{�S��g2\�m�G���� �t�R�v�"���.���p�Q���zN�B�z��!U���M���ڦJ��l�d�0�6'ٛ��x�,!�]���*��n;��a�=~0��y�w�DMa����xC�C����O�&^a�\�r �X�`�+�m� �dGP�'��ic�z�
Y�f���Î�34����+j! ӫ�\� (���z��ư30l� ��F�\�s���t��H�Â��f��_�������~WϯZ�lnɅ�Z�z�	�k��+��g4m�~*d�����3�<)=����%���qB[e�E�i�,��ʭ���{��i�|����x-ē��[k{w|�%�7Vc���U�v��QS�ګ�v,h�m�T������є)��cުw�C==���A�b����?��N��$d���u��s�v
X�6`^�3`6[�lp2��,�9�����kh�: l��^t�=�1u�w6uw�*jo�7z��ʚ2e�`]���mÎ	z�#P�2�Kl�;Wb��5a�7qa �;e��c��x1�v��n���r�AZY9c�^ߠb�������.��j�z������h��5��B���@8�����[2	�p�7�xW����t�3��dY���n��|�pO�������:	�^�	Cz!6}M����Gb�[�җ�
����������ޖ�{�{�f�~��>1C8Y�V�m4�IjK�I�ĳ�����m�x��/,@�M+�i�r��y�� ˜!��6b���g�p��3�#�Q<_�y6�\6��k�9މ������"�1?Y� ���yD���~Rq�"��gB5��`9X��2�@30�
O�1+-�5`L�^��B��Ya�X�W�z`�@�X(א��A�q��j��B�G--%m�C�
�%��_Tk�=�h�N�w��:��6� a�{���-�� ;�)F|n��q`/��13Jjz1�qrRr,� ?�	���o��1��� �e���L�8���[ߺ��4�|�Y}�+�%�|����/t�;NPw����W�>A�W�k�z��q�_X8�r��y�>��Ǝ9�c��U �f���F�����-��]�q�٤Ћn�1�@��;�I&;�:xŏ�׸�QL|��u�]7�g̑�6>"��5)[&h� �!}lZ(��8o��6Q�v�*fet� �n�]�C�>f̎�2�����ư�gN�I�A�����ߣ�v��c�?D�'��W��%%�q����*��� �p�ys�־�NW~+@��:�	����)1hDS~����7�12�j�1&�+��gZ���u�1�t����X&���Z��}�/�V*�������9��R�K�B�~��r���g5c�#��v{�^o��J�.��pZ)j<&�s&f�7h��Ldg�6�ۺm�p?P��8��Ƅ���B62��z0���]����F�]w�y? �㫥#�1;&Wj�c�=��8�<V�8��t&[*���3��}�N*O�6���1U�����S�A�v 뵒�}��Q_�����t�E�PlҳOm�ɧ�'��Y��Xb�[�^���:{[��e���Id���v_L3�X�̴=F���Gh����J��h�����C��بZO�γ��T�q���;��Wb���K�<���z���;5eJN�~�l�r�q*�K�����>v��Փ�G?z�f�<T�2R� 5�pO� �d�v����������Ƅ�ޞ�c5�r�5evmF�8�1�އÞ��S�����n�a���O�x~q{�/�0g���#��bU=9,�Vāp�q+F�:;ǒ� �w�xq΂��f oK���ټ�L�85 ��1~���V�ʽ������k��L�?|�cz�k_��˻4��w��/�Z8�4�rν�[.~iFb�ܰ1����w�(��!��x�c`��bO����Г�x��	$6��+1����Oa�e����x^��X�����4����X�z�]��٧���ޣ���v�5i��iμ��S�u�~B?���i��]4���{����2A��^g�_�<,5�qK�����):�T33]�nM@Lr�W/��egP������+^5��>�ûW�/��2��|�n���X�%sj���x���'�yaq[����ld�����+�����]c�Ke`J�Y��mS��O+v4������|f�EV�~q�>��k�裿R�(}��u��k��>���3T�4��9r��	N�7ڼ�5�@��̀��`�El�����ld����D����X��(9��]CV��Ɔ�-v�F!fk���EX?ӆ#V�4��;^��3#{Kq�ʆ����3���I��x��A�Y�����8�kƽ���i_3;��`{,c���X���G��sZ�d���vU�]�0��_v�N�}�:6v���\���
m��>��ŗ�W��-iܸ� �l�pQw�0;x��զ�U���Fh�~m���Id�\{%�����#BRvt�m�.�4�7wЇ��wY�Vΐ ��|����{��K^�G�_{﻽��Wk���ԓ���i���R? \�	�dan3JY����q�B�Vi��̛,T���꘻��1���d�=��1�1�z�!FݴR�3��Y|<��p���%6i#3��6ǋ7i���5����-�L�c�g�n����ux��������Põ'f���G[z����%��J����t���ּ�NPWW�>��O�ޯ=��^���ϿR{�}@8���4N� $AMn�W��u���A�����i����:�����%�S��M���'��^:�o8�jaœ4�vK���{�b���S̄c dW�po�.��|��kt�st��ǫPl����Yg_���A�>m&<��s� 3A�v�?n3���bOz����eo�@i���ǆi�g 6%��@�`�4;����wm,�GiZ/�&����u�q��:.���ٰ�š����H��c���4�r׻<"m�Y����f�Eǲ�Y��ѭ�W#ݗ�OCK�-��E�T�/������Ь�oP>W��zH���۵�#��|讀1�p�Q�?���4��$���s��z�`�n$|����0�Ɵ�=��0؀f���&��f��N�'�[��:9�Տ;�g�Q�qU�+aO������~��ϴ��4󀝕-t�l�������Q�:Y��,���ԱH���1� �l>�<.�9�k�� b��y���n=��o�(bvf٥�ᦔ5f�1�ĉ��i��������b&2T;�No�u��Y�~Y�}y="�$�%RiO��c٧��,6�d�I�e������D��!3����1��Z�sҞdl��bj[<��� �|ų����]Մ�y]qջ��YGhܸ�J��V���������M���z{)yYT6_V�ZQ��2�$�K_�� � l����H�X�{�P���5��_�翢 ���r��ń�pD�CVʴ0��ck���1����Daa��V�� \��Զ۶i�]�iC�RU���6^O=�^�x�ձ����/�0�-��>�p��@L|( 5Xx"yU��{贗X>�Ryp���'!���s��k�a?s�v��4��[����e���������:o����>�}�����C�q�؀�k�f�#M����^����Z>������>���Ǜ�x�J���,3��3����� �ٚ��x6�`�Y����>��$E-_(�T�	�w���=ڰ��9Wrr�1���#Y)S+)��6�H�9ֵ�H�H���M��Ga6kLY�zq[����@��t�l�(�$i �d�=#	j���<610��M�tJ�����U���d��Śr�>���[�yd�>��E�x�z��ԏhd5w��6mor��c��L�>�x�P�|S���p���"fαu
�Gb��.i���ń3��3hx �gg`����(1�1�4����)�!p��2`{\b6��}p8Ǚ9��a�5�vJ�A�v �Ά�����:�a挌Y�w���<֩��7��/�W��'�I΅���4i�8͝������Z�̙J�) oK�d��m�f�LQS���J���`��{ｃ�ͦ͞�B�)�wsI�����ޡ�<_w�u�t�Acw�\r�|z��FCeGp�=B�W���c�.���IY<!͔�(����Rw������a�������h�굡�i>WRSsQM-mZ�zcP�z��l]n�5wΙ�6}/re)�	dN_E-f/���7{��pb���}��J3]?�{CM�l}�(i��B�H(Ļ�x�����c���H�����H�7���oo5EnT�Q�:v7�vV���En0v ���N)C�.��i��R@�<Q��=���cEǸ�]����x`���Q����Cޜ�g\�ߴ��
��g�����/*��e�i����	7�b��PO���,5*�8��bSC��^�s�j�U-��:�����k�T���G��H�.��L(?��J���P�O�k��M�{S >�}t�s��B���	Xx�x���E����\6�"@t    IDAT �< .9�03-����SY�z��.yF]��SsSC}}��+W4q�d��Sn���
R�0�����~e�y L��2��� �!�%Č(�$b�|c@
h,���D�aƘ]��9f�~����� "��ras���K��ٟ�/n k�a!ŏ����8�m��|츞�r?p@���� %bx�Ϻݱ��?:D�U =�x�ϊNS��
8s���T���=��C������9I�q�Ɗ���U��<����̌�p��b8oh,w�g% �U�G�r_+��^ݠ��L�I[��TTSk���k5QV��ZhVo/ۍ��q�^�t8�ۃ1>>�}86����M��?��I�qɺ����@8��|���ߘ2a��<��([��B�0���I9A��A�cX
�,�5NQ<��}�׊D�< L^��{�A0����MM	&ŭb���[�1P��(�ٷީ���ڸ�O�Ţ
�R-�\�k\���ԝN��>���S�<R=a�>���A���4x[�.��Z�(iV�sm �ﲑ�Ԅ�a�Y�}1���s�x> F�*��� |�nP��ǹ_���:����� � ���\Y�y�S-p�sJR ���͐�5�w��FJa*ڈs�1l�g��ϸ����������h���Av(�� ������ (T�s"0流��G���m=�n��A3=��3!E����^eգr��9�/kVo_C��O�{�|s�j���M}�l�h�:�3#����/�)�<m���m`��L�^`���p�=2�Tb�|"	��=�^'��z��#�q���4PO���^{�؂���~h�Wߙ�XHKk�jՆ��ݣF��LN�����S�冝�1�E-BA��ꔫ�4%��A�if�Ii��I���B��̘1#��b ����G�v��@>_U�����[]{B�x�����>Y�>�<��7�I9�F1	GL�'�!&A�ˑ@0�2������l �FG�A)��Åtb�3[��5�$	�1�iv�{�:�|���L$�0��z�{ܟx�ĕ������R|�S�gr�����< 퀅`L0t�{�Q��Xo����C��<z	�@��u�6�S ��)�އz(lЁ���^@Ma�C�e��w�>���;E���.^�zU�����Q��K;m?NMM5��!&\�6i��u��ў�LW�RV�*e�.Ԝ
�$�P�` t/��2��#��b�9c@�c\���!��˸!_��(Rp=0�3���f�:��y�K�w#�����W_}��u��#�Lza٢���C�[���+�3�X����*j{�fO|�!m���Aa�f`e�H�d��Ը�>��;�4����5��E8������B���/|!���$�bya�@d��Z@�)_R��1�1ǙX�b5��<��]r�U��ͪJ��=X�=�1����ܟ� \��u�Pc����,���3��k��r�,>��y�G��	3�6�����0^�������� ,�8��(������\�������N1�0
�t�	0ia�0�ab9��w0�i���|Ǆg�>����y>���  @9 ���+���Q�T^�I��6��x �@tC»!����4�q�Y���[�C��p��O=�{�v�*}M�Ь�Ν�N<R���pe.ӦR�E����o_(��VON�A/���`��?��3/��<)g��7�9��c]5/��60Y�������1cl�27T=a��������{ǫ���l@���\sͅc
�3ϻt��/�\4�^9�R-)�ɫ�WSKKs �=�z��>������lM��lN�q>�7��(��Q� 1
- JO=arsY�Eh��T����[B�O������}3��,ۮ���T�8�+���o���M����i���R�@��Cج1�lM�w?�s0��A�ﵑ`���i �;� f��p^��ű������8��V�,�@76ʐ��bHc��Hߨhq��k]q���' $��K��γ�O�-z�'N��st�I�u���Ћ@��v�Oȋv�=��a��-�����29ai > ��_�@�0l�5,��q0��C���v���^r���0
��c�6Ң�Xo���z���s�"u��P{kNW]�>�=��z±�-�m��ڲ�{Z��YW&۬j� :l��K��.�{���M7�<��|�;�O<��`h���y��o�G���u�܏9�0n�/޸��r5�r<�x������"G�����n�馋��o��["�M֎ ��ٰzQ[����R���&���N����4Y�Oy���v=��s���,9�f}�a���Ą�pf��~����N�q,��p�
��<(?J}�y�k�UB�?�Ov,k�<x��y�Vؘ�e35U�6��?���ݮIo��Mݶ5���S�:�̋�ݕS�)�� ��i���*�bx1����
�X�Ǳ\�t�i��q
�9�Q^�H�2R8"�	�����@p&Ɵ~�)����7s�<��\ȡxU +z���5��	��q�y}���C(��`�.��;B��"��<���c��0�	`��:>G/��LpXυu����0fX/s���,��9j<��Ah�?!�{ˑ���� �乧�h�������Iͺ��s��YG����J����f�~q�㚶�Q�i��jd
�د����F������#dƸ^q���Qo�8�s�!��NcG� ���z��y�������8��$���{�a;�������Qq�8 ���~��7`LAxƅ�Mya�����'\)�B)���6���t��o�#�TO>�t��^f�h�]U��R� E�����s0��8��f�p.'fP�߼����x?����)[�8~�������Ї�SO�
�9�x}��sU(4�G�i�T)����0y��%������B�����p��V�����E0*�a�L���c�~�A�r�ӻ�Frg��c�n&LȀ��SB7ƞ� K�i�f�q̍�1	a,��3 {�9��yc ��|H� ����[�c��41���]E���B?�D�k�m������� x'c�w��ť��0n�H���n�ﳑz% vs��x>=��i�s�W��թ�m� �s��Je�~���u��Q�:Q��M:����y@�Y�������R�$��	��� )tQQ:� R�@B�Q�qG�QGfH�
�{g�5�;cEE�����S�~�o��9��rJN`֝�u���[���{?�����u����!G%�R��e���S��e�]�!8�b�40S�Pa���I�A��ڬ�3p}m����@�/�'�6�ߋ���q�8+�J9��>z�=�\7� <nժǫt,��nڬ�u-:����w�Y��z����ٙl�G͆��X�3o�#$�iӂ`~����b
6�Z�`��0ر�! ��1U𽽬�ۢ0p���U)���5���1=����k�F}�>�IS�虧������0�#*�L��-i��Q�'�[e�=�A���o@�
m0�s��km��@�s�n���¶����{2pa~ L�Ś�0��L �Qz}�*�E?-'�況P�3A�����Y�q�#��JPl��͎K<9ޡS.�ͽm��;~g��Y�@p/ƻ��k:r�c���B6��g�s�"��+���e ̭�������K�葇����ujn,k���u�Egk��պ��껏=���?X�}t��r�r� ?t	iJb�y�<�@_��W��6p�g١���?2¼ cb@���l����y7���#ք�X��i����X�ڛc�{�k9�N�:u���Y�|̠������?�е�X���">�g�q���6U?��h���P��0����a8��cDg�Y�`2��.x���E0<�C�0@�{X�:���zo��jG`��li���;tӍ�ʕ������go�[�v������U�U������9������Y7xt�A1��	���OWA��L�׈A86G����x�̭��`7Р�	�g�s,� 6MLV��@�Ƶ�m~q�P�ν���ڒ�	/�q&��;6�p?�1cԑ���dd3�ׄ����9���Q�C/�\�~9���v	 �N{��X��皱���s+C-�C��+��+_�??�U�^���h�7|Pg���ڸ~�n�y�~�����u��kn�aG�R�$�K-�F%�s�r����!?daYǋ-���6;X</��wh�<�gd�Yg�ٓE�9���>Y��+��3���g��= �i���	L8��<r��wlXA���u+LLW���� ��艺����Ц���7!D�d���6?X@�$ L��A�N��P�PW��>еM�	�c;jB���>X��dprj*��#�*��<h��C��RG��ϿI�-�������Kws��v�<�
��Qԝ���t��P%j{KY���0�OD&p���A�,�����bu���|��!е��&llN1��J��6�x������`WM
$9����`���C�T��Y��ǹ����E���W�C�`��_	g�K�����s�Ǝ�n�s�{���U��/�;���Ə?P��Z���jsg���Ň��(���15<���}�� �L/�>�&*k���b�.����p���P��oN��^`?��o`�&���D�Y.�[�VK�l��;��������l�w&:b�����sgiźez�O�14 t\�դ�	 �ax���N
�;2o̚=�	%���k�q���� fT�/���V��t��1gGV�a�WJ*tm֜[?�be��=�T}��3B&Вڃc� ��l����9"��3��cbS��3���O
��|��a`��8���06ؔW�X�1P6Ma�m��?@4`1��ǚi��_��@����w�cb��5�Ʀ����#��tQ��;��+�e�Wj��_W�k��[*�w���5�=*:���	����В%4�_k�}�W.�U��{�|�a��::��
���%�\4.�M�Ih�?��OA1`� D�s�	6\L���ڷA�"䎨�X3�0�e,d����R.���]w�qð��W�t��+��7Wߐs's�N;�T=���kɲ�!l��au�����@��`�ǃ@ '�pBx(؃Kj�4;c�Z=��c����q�Οv�i��.��%�os���-���ҟ�����cu�Q����|OIK_�Ѭs�VG���%�)͜y~a�\���µ c 4����w��?1Ǫ��A�ks/<Vsm�����LX���ju�{8���; �m��N�Ys/�^�G�5���s{�����ׂ�`�>>vG��ζ��8��h�zh��
ɦ�7�tipp74���Ӛ��z�wK��>G��q��ne�Ⱥ���T)�T*&Yq؄!bk^x�L!bD�xnجd�/�;�gy�[���0W��=�v�����0�
3' �{�89�lF���6�';1W��b6���Mw�����&L�ܸ�5��[�'c�舷�&�z������֮_�j�B�b	:wG��xP�^1G�[�����(���
��*��w�}a�
D���g�\/o�9"�x"�S%�/k:M���&˛5z�D���M������`�% L=a2��L��]�]���� �An�!FFqh�@��L��l��M��`�Vk�����^`��MO��$f�Cɥ�����5�m�����p?�9�K�J�ٶ]y���z�٧þp�Bݕ�s���Y�P���U�~��ܬ���^�ƾ.��\����A!�����&-��5���D��BRc��m�D�x<:[��v�����2�L ��	���1�W,���}cre�nظ��rJ��o�}��ӦM�8�P;b�K���g����<��t��g�W��^Z�2�1ǖ���A���#�!�=8Z�.���Y���r�uׅ����}�J��(�m���/�� ��@�-�m_�p�Gi��mzy���Ve2y54)0��Ͼ����_�ё؂�a�C'k���>fr��D� ������13u��P�C�p��X5�Y�ꟁq��
���MW����Ү��L*;bnٕm|-�m^�jY�Z*t��Tt�������fHDO�(��yO55�r�.)ϙ��A!���=}�����`�2����n"�K�1cF0;����{��̙�����:����;�@-��B�YͿy^r<� �p9��磏>����t���΄]E���9��դ5���4s����y=�̟Ö�v��c�p��!AN�Dh��@�`��}p���#,�3+S�Y�3��6�$��1 �U�]:SQ�5������6mH���*��qcv�K/��Z��v3��؄��>s�4�J�ⳳ�~zU��E���t�9��[˫?�i��sG 8�����֪ݖG-�0��YR�:_&�� �Kj��4�������l��*vwh���ҩN)UPW���B��1z�)gj̘�T�Шb1�J)q�Y�1�ݖ�3���μ�|@dy����GG�ܘC�B2'a�c5q �դ��O�+r>�&�{�������.��JB��j���w]���V�؄x�~:��)�(����R��x���6���z�bV���P�6G�9���{:Kܟc�<�b/?̖�!(�:�q��*�h�吨x2yңN��CJj9�wu�I�L�:�Ⱦk�a"��:w�y�<���A �)q�ݸw���1�:��H��;�m~qm�y��1���w��A#��Im;�N�u0������<�%��xQL���j,���ᯠ���W.��a�L�	���\���TW?N�BZ4I�'�|1qd��5&s��^s��z��fln�{�Ø�$1K� ���;���!a�1А�B}��_��0V1� -����&#'�6�J'�!j�̷�c�Ǐ<��u;����-���=E�6jB�	�a���o~��M��c@@x8� ?�,�4�,��:�<~#�{�w��� ���Q3D�I	�A��2��y��8�!���,:�&��B�[�<��
��rlwTج�&���kR���p5�J*���,��w��D���88� b��<f��q�c/���1�m/H�2P˯���}����<����As!��ׄ�ϵ��U�Ȅ������3=�yf�����`���x��C�U�$@K��|!�l�I�N��Ɔ&�����T	W��E�x,|mj8I֠��F�4,�^��l3Z���`8�v���a�0a��!m�9���F��m�Z8!�d��l.�J�\6��=��9���W���4�	7�7��Q�q��3��G+^Z�%/,U{{bǵJl�<�l5��WNm�{-�f5C����k�C���W_�C9��%��	� ݡ-�U���1�[l��Bq�~�����I��Sg��~C�ʩ�ҙ\���3�Sʒ*jea�I����L��sF$�jI��dj�X�g�v��;锖�\�i=���w�j��G+�KJS��U�u�m�}u�1o�GLS{GQ�JJ)�WJ��i��������R��K/�4�p�l�/�	��~!H�9��)���p�{�w(h���66�Ӭ�cC&t�����ߞ;w�u��c��qkV?4���V*�:d�)�������8I�M���Ͻ�ի��q �M ����0`�}̪��V�">���������b��
�*F!l4_��8;�͌�cε���*}:C���*�4zt�Ң�h�2���x���o�jU��� ���0�r��3�Wk��gD�!�W
�.Z�@ULu]~��q�)j�˨��H�Ѫ���^Q*3Fi�V��R%ӭ\:6�����Ct��E4�B�3gN��w�D�>�8߉~ ��sX  c�.�1_��`Ä��DJ���t��Cr�Y2f�6>B    IDAT&��];Y���R��调�����	Kt;k���!��}g���l�֭��}6^Yl�WV= ����P������v�|�PҎ)�1o޼p�PGTH{��߮�|�3!J"V�$f�-Ղ���L���l�F�ɨ��U��l&=��պ䒏�u;4�
��JF�g��)��1W�R�`����pL��k�H`WH����5�������h�u=�3�ÚuJA�,�њ�Z��G�R�Z�^�|-2�����K�Z�,;����>��`������ʃ=���������!`�kӣ͛�/����Ô�(�
^8�ӱ���W 8x��_�"�@�l`�Zeg�]»mX�P�uô�� 8i��V�iJ�I���ScƌN2�÷s���8�֋3&U{,3�_�g�(�DG �ޙ��B��te�`����C�j����L�ݖ7nX�_��:���:��7)�Mj��y�K���Zs��E�% ��1�P�	�����
d��&�W
����}�+�fRjn,覛/���:Y�9�TI뷿y^�<�J|�&N<P�JS�쳱�.D�
�`I�� # �@|�C�8̊��d�'����)TX�.	 g�9��q��sc �?������kሃ0�&*�Q�;�7�R�T`Ι3��ag�ׯ[Tױ��Α��-�C=�jW(�<��#t�'�% H�H-�l���#�P�����s�y�sQ#0�� ���:��x�� a��Pq@s�6��� �J��u�LݫB��>K�&�Ջ���}g~@�B�*���� 3f^��p�3�g�`^�WmF��hD;(�W
�+V,�c�������-��NU:UԿ������Y�^���O��1ǿ9�
W*�����F�f��0�ǹ;b��Թs熞�9����.�x����M� �DcqVᓊ��#ށ����)�@���E��.�qkW/_-�@�#BԚ٪VTH��DB�:��nq��,�S�(BA�t���PT��8�թ�t��2樂d�`�5]@���  �`&�ӏ���s6��hR�ahwΟ�g���&�у��}��[�?�R]xUH֠�O(����3߯)S�Y�M��F@xg����m$�J@���M�ڵ�ScG�t���k��wjs�z͞s�~�K�P��n��Nt�a�(�\}���d��#�a�c��Z�X���wp�S$����q�|r�q0���D(>;m[1����ua��;�Zda��*�e��4�8[N�ӏ͝;��ag�J�
�`��$麥LA��u���ӓlX�-gX�xKE`�-� /�W�w ��~��E�Q�ױz@�v�@¶'ՕԸ�w�������	g��ޭٷܨ^���������c�ЦMy����U.7�,*>�͜y��L9<DRT*���8i��H��p�@��RwG^������Ӧi�����Mw�W��V��s���a�&M>\)j:gɈM���٤�3�"E�Al64��.�|��7�u���8��q�`��7{�p�5Ny�k<�b�`Q����WųV�Ȱt:��.��7�[�n�xbsKc`��1WW�Ls�8��)D@.�B����u��Q�K:㒌��p�w�:�Շ��pC�\[4Ǻ+��&��j�^&�V9ߣٷ^��a��^���M:�Ѓ�l��:��K��7&�,��`��9+1G���4��3S��.x� ����z���RW;󮬹�]��3OQ�{���>}sѯ��}&��+����NRO1��!	_���͈�\a�q���\O��;v��������l��̆�̵��qDD���Ys<��,�h�kJD �zX�����V.j)t��ڹ���	��	������$����N���d������w�WBg��0O�	���3��.�|����k5��k��tj�y�ꃗ����F=��5��k��ѨR�Q)�Bh͌Y�4y2;�ĖOU4�W�17��C�8֫���7*����.��9fq�
�0��5TD�p��p�^�&Z��uX��q�'Em��c�]��>�~��,�=m����N����R�O���~���};�;`�y���qV����{�BZ�u[MB�w��0��'�Sr�!r��Mrh�N[7PL8�6����΂0��d�Z�`�J��ru]�u��������e=����_��^x�U�l��v���^�^9�;���/�����1i��L-���1N5�|l�O�����׋�.Z�ݖ������]�vQK���0��qN����������5�<p��W2l>0aq�m�����3��!��I����qi��vh��]�������Q�JS(>M�f̚��p�'��T+u���A�=q��n�\�Zu)��S��"��p��<�'iF�G�h�������l�LV�8�k�-�1=��Xc��xΈ��#���/0n?�f�p�'�.��@j������g��}�N���~�M�+m����<�6�ݬ*ŋ���ŋB�:�+Axي%!v�T(i�>y�L�q扪���֤��m֓O���_����J�:��C!����I����W��W��ߛT��oG@ئQ����\y��NL,�g��wo���+�u����X��'Z �>�@q�H��^f�NQ68 L��	q��y˽0it����=V�2��mVS�h-{�]g�y���f�������A��)+�)�*L���꓋ۛ�=F�q��/���;9�s=x���:��LĬ$vV8����w��^f���t𻁆�9�����r?��+m�6��?�q^L�P�=Z�4�\����̺�6G���g�jp��o�1�������Ƞͽ}_��>�{�c݋���0ǹ��e����scW��eID���.�4K��r�f��N54�U*d��쮍Kjo/�P��u!A#��͙�b���W��7_���gm<������ZY� cW̼��S�����+�9�U��|�Ec��'_��v_�jѨB�I1a�[8�zŝ��TK���|_���\fC��9�7��p|ߪz��vi�j�H�bSV�j^�BU+���K�/����*U3J��	�8W���5�����d��3�����d�i��'�A����,��!+&���kX����f��z�5�̽�Um���l��p��f}6�����m4�Ƌ���'&��^n69X}�/N����	䁺o3��������`��˱6�Y�f��a�bD�bY[�q����V�I�A�>�Mܖ�����#���bL�Au�4~L�.��]z�U�E�D�R��S}ݨ��y}]������f�&c�d,Jxq��3��qw�ׂv-��u��{o[�?��+vc�Hᜪ�	ׂp̸̰�[���9H�����ʃ�5h��vA ٢�c�~���Ժ5k(�r��r�z�*�S�ohQ)UV*]PEe�
�#�-���(��ʹ�K�<�'񍞔V�a� �����4�&����ӓ�L$��a�-j5׌ˏ��!k�~�y��<d0λ7��b�N�`�um�6�Ӷt����ك\�u���݋�˪���=��1+�6��5G�HUl��d��W;��3}����!O|�u1]��y�~�����k^di�Uk�(l��UL~�?��GWV-�hۨt�]�P;K�6n���{�Oz�v�c/e�.�N��t�Du�)�6���M��˹�������cR�������~@��y�Wu�Q/�H[���c�K[
�0�~A�6�n,>��b���U�xL��~haN�r����sO������IM���F�lV�RU��8�U@�"M����[� ��;k��h3��K�l��$�0Q)��>1	*�!A�	j(a7Ȉ8I�'��_(t�9 $��Z�����'� �qA���d�=U�l��b�]p�N��dbq0x�:��ɉ�Ǝ?ˀ�L~��K6��L{�;X�Z��j=�|Iq �+�^C��I�B;�XDlF�:�[& Km�h�F�i��XB&�.���m�t��yCO��g �\YA&X$y�ĭ"/�̟Y6ϖg��[�ߕ LQ��}�U�lST%^2!r�v��봹�K�:Y�l�r�d�qU*�{���	O��Z��s�x����rCͧ�߇2G��%[1h���]½���΂��
k üϷ����b��̭?&�C%�7[/�淿P��LU�Rw�l�ʤ���5&@�) <�d��a&7���%�� �~3��8��p���0)@��JR 79�8a|��\yw�1�9 ��K� �g�@1񩻊�)�xҖ_���xF�-���m���B �v�`��I��Oo[*Ϙ
ZLt�B�8��}�%�˽�~�\3��~�0� ����CF�G[��"O�I�*�����!��ܗPo��bĽ� M���:,X,T���; ̋E���vȀ?τk"K@��Bv$, /G}�4�+Ax��������J^jl�W�ܦ��M�$ �󅂪鴎<��e��ZM�.���WM5�.y�8d\ׂ�@�n{�����������= <��ˇ�9�Q�)&<��QadC��b����1� �؛��\�kS�j��?�C֭U�ܥ|E�[�M�ղe��kV����J �`���c�2Ø(v%� l�	 ;X�?�,3�aF|���9�&�yp<���
�	l  P� HS^�: nP@���H6��`��I�
�'���Yک���Ϲ ��u�v��~��<ٶy �̖{q-&�h3��Q�q�S�C�],, ��� <��*,<��s/��>Բ939�Ŏ�xN�'σg�,���^ 8l�c i�N_YHXmd�,���`[6�;���b��<{�gjA��^�M����c�}G�.JS�5����&�^T�浹s��~��z�[߭}�>T��U��3���9v�B��l���V���s{M��.B55��Z3���]f&Nx��+5�;O��φd�TgC&$k�����r���<B1(���*n��U:۴�X�G��"����L$۸��Ô��;?<��L�#�>w�)�U���ՓߨƦ������*��Z������Y��z0G�5�bM:�e2d�kA��2�`c�!�~� �l�]�:1��<��L~ؔ��Ӏ�1��<X[G��#�r<�@�8����y����� X�B#{���\� �xN��H�7���q.ㄾ��{����?m`���������S�9`gq��� +�8�|0K(�A.Ț�T�b���A���� �bd�����>g���g��u�xq��;��MH ?�ݶS�a!`Npm�X�I�,c��{7�\�bqp�mZߪ�v��}�l���ǩ���r�G�ι1ڼ9�je���VWwYM�Yu�t�:�����Q���Qf�|�]܋��X,s�`<ύC�)��e����������No�����4�|Otļy����/���ܴza}��̦Hs}5����P���Jp��q��OT�J��{6�L
ob���*��t�Վ������d@�v����������	�Þs�r�z��Z��S]t������^
;̚	���Fv�M� l0 &�6��H>��C��N�(X-�������W�@� ��f���0���G����C��^`ŨͰQ��8R���X8�@���� �˱�����xؓ�aV�7�����X!;=c �9�1ǀ H�1o�BΜ���&���ڮ%���{ ��XlXt�&�&�"�<Y� T�@�]a�L��&���dK�i}@saQ�"_�c¶g�"���ۆx��$ WՒ�/�-Rg[�Ǝ�j�͗�BX�t�ڻ�4n���v�mzmr��Z���U�b�++��w[6C��k��2 �w �,���f���LМ�#憝��a�&*�D�d��D���`G��J%��'|հ�0{��~���ζ��)�TQ��O1�W]CN�<�+%*��� ��#<Ջ��g�B7�5x۩��v�#`;U�jq��"�@�d��!?y�3n�~���j��M�[�:M'��`Vk�t�S�	��JՆ�w���5�� L�"|wu5;��	�2�=� A����dE^  �= fnL| &� 7&7�s`��x��+0cB0�`�� ���po�wHh�L��6/ �q�[�\a�,V�9���l_f�� Ф/����-Σ=��x�^��π0� g�q]Tz��
� ʹ�``�˸����3y.��p��EF�l����2d� [�s.L��3��3�9�;r䙳��o��bf*}�0h�:Ni��%z��_S�R���Ҝ9�駟�;�T����	=��K:d�������Ss�u�t(WGQ�d�O����5s5˷&l<�fc6���M��/�\kb��	��$yZ�&��e�}�	1G��r%��~��{����-�w_�baK���lu"@�R)+�n���'L�-�؀R�H�B�L�o��V{��v��F�� �J8�Sb�39 ہc/*�������)�Թy�����6o^���G���7d��S����_����JҖq(�% <� er�����Ң � Z��3Fd�V@��
�,lK�X�C^PX2e�H��°sO3E �g �ƦG� 610�l�@��!6Q �k���}��2 3�M�8�>9��`˽�D�%@� sM��Eơh��1���P��	�v���B;+���`��]@��J�3����"�2�9y�Ŏ6�Ok�Ȝ��\�5�d��	�̐?��5h� ���y^���?�+�l�KAx�KZ��UK�Jk��Ϳ\�{�z���ӟ�J�7��|OVW^s��8�DeӣT�H�2�T({03���GN��y�hO�ƳD�@V��ĵh<_�<�d��r��q<���D�geG'��:���W*�
Lx�A���n8d��Uǔ�Ǳ�Z!_
�,)��^h|��@M�vb�`GC�\<�a	�AD�a��n�4�z�:������78T�������N;P���f�m<n��ݺ������뀃���7�z���/�×~Lmm�p�Rզ^&|^ �lu
�}v~��&��ʢ�בpV�@�LP~�%�¶+d�JS�=�vu_�l��0��'��sڬ�c��)���ن�p��{  fl<&�:�~�xb0������ar�x�~ Q�f��G����1�Vo���N{i��/:|v�/�O{��H�s�#m������<g��$�����lwx�e�}�䲘�f�5�v����ыK�롅U,nV}]�����f�|�6ml�=wߧ�}�7�m�7�7ݮI�O�]=��R��d�Ą�{ĝv�i����(������a�4.>Ƹ����7� [s�Y�vf�c�@:x�g��&�q�K���{A��ٳgo)K@xb뺅�]m�3�\�	
y������+�q�����eU�����gM�`m04'��@C�`��j�đ�n���\F����g6��Y�A���C~%�|gE�n�E�?�+e�6����[O~��-[����a�{T��$LX͚u�&M:X�\W������=�j7�b�۔c�*�M0�����;	��������68��N�>������v73�Ë���+,3:O�x�q�l~�M��VK�����;'��teU���Y�q�9����30����m��2��W����Am �Z �Uf'����8b����8(�}6�N��6~w�`����#vx�c�˖�������o��	ҭ����N;I�m��9����T��{����M=�(�yerITQ�i�*j�02@���;�`*��8ϕ�Ȍ� ���������52��*�k��XC�q��@��,�D�`�w�5��s��t��a�Y㈫n:t�+d�[��A�!�uww��o�K���m����i���a(m�ST�Xږ��6ͣcѓ� � �O�l��7T9>�+_	v�3�8#�!��F������ǜ��+OG�    IDAT�+ ��ڭO}j���ԏ4i�x��wh����3O��%L���T�և*j��9��!�vN��.6G�m��N�X��@��6{d��r��"��;�œ��s�rA~�4l����s�����3�y&#���ʽ ,��g���|���Ά3�X��Ȃ����U_&�ߛM�U#{�9�?�JdO>�iƖ��N!�B�9����=�!��Ym�4r��zA�>������{YC�Y���SZ�b���Ejoۨ��Nͻ�]p�iڴa�>�/�_�ן�Ҳ����'t�qǆ"�
�d[#�Q�p�9��o���l�v�7�g��}.�5o��0v�����O�<L, ෾����*X���8��X���q�E8"�x���[���r&�}��9w��i�h�G�Z�`�JǱ�g�������t��S��w���Z&(����O���)�L�1���c�;�ٝY	��mo{[��~�{�9`G������������I�A�9��=�R��n�2�c��X�]v�>r�tuw�h��]p�uj�{[M�#f]lI$v�����Q�X�/��<t����'��fu� n���,/��|�sl*�y�A��s4��e�@����ф.d��	�1b0�������@;=�j�7�r���%���k�6��k��rl�����w�s����}N��5,��vm�#�ux�ŋ[��A:�%K^5���E�4�u�-�j�̓�M���_?�O��`�,��Oܦ�'��ik:$h�v�9���S5��1g:V�BB>>�<�����*����
��9�6f������9�@�߇gRL�e��t��;�뺩S�&����4m�L���������:{��Gu��}�;C��~��:;��
�xŬ�3 pf��`KF��>�h`��G��X_�@�%�53 �=�s-<�cV���chS�"���z�ձZ�<�kM:dM:l/��}�z������nVkkZ�*{�I���2:k�E�t(E�]E�]�� ���<�v>���F$�J ᪖�X����ʥ�V���C:�ijl��:�z��.=�41�j�}Qk[���L����جb>1���	���}����H,,���4l�̗���}�-� #�r���hD��W���	<6=،�Eڡh^^4@�4m|S�F'�(���J�J�\��;����
�؄'��]P��z<!j�i�6��N�!S������/�PHV�����%�ۅp<������?6�X��a' �����9�;Ǹ���5����إ����R�s����ܨr�S�GM�_�ިY��PwWV�j�7��f��v|��Z�gϬ��tF����.k��%z��QCz�T�М����oR]}^�tFݝK��W:�"�T�dT�P��v�b���0G`jt$��ؽ���`���7�	0��a��=*�^1{bv�s�5�X��и!�6E�u6h����������RK�l�����#�<rݎ�A�0 <�u͂����c��e�5�y�>��KTɕ�_��Ouw�H<��Vt�^fb���x1n�i�Y��P� gױ���TΪ��w�3���� #�4�#x��n˱3����nuu�V�ؖ�vR$k�U*JK�n�}�}]�6��	�>��532G`~�-�/T�1�����#Ǿ�0���/z����zM��%}����䓧�P���J���,��'�\Ɇ��L�M<��3qj�",�M{�ñ_�)�NҲ�Λ'{/��$�g��@�W��::�� q�|��l�	�����a&���OÄB���e�5o�m�s�1�w�Y	�c7�Z0��}<�ly����^�v�~�įU�%�/Q�a�?²��6A��*d����'}�8<�
v�����á�V'�Թ'������ Y�X��?�ca`Q�uVUPO~�~��k�3�UW�S6�l�Ġ��(�kR�C��I�U6�c;�R|;"x��@����;z��G$�+%`^��y-\�U�Mj۸I���'�|s���+956NдN�!�r%qВ�L)K�r�]3��π���K�%`i���Q4` ����7���XjL�\I�s�CS�l�4��\���8�,<�`|�;�	�'LX�\.�y�n�İ���+>y0��K=�I�8���u�Y�ӟ�{R/,Y6��� &:���!^]Tg� l������P; n:H��?:(������Fx\�$�jbo:�?Ɋ�.E=���*tC��J�;ܷГR:ۨR9�ԎH'�`�	;:"��� �����n���~WN��k�H`g$`~a�sZ�`�*��+$tmV�ԡ�F���PS���>5z|ؓ�2���$�48�z��8��sDQNl� N0�a�~�l'�v����û����\Nہ�>9d]:���o;|a���G`
\��.��A�j�C1��,�3��O+��<q͚���]Ӽ���'�E�z�;�ğ���V�8�L&�c_1�I�\���Kh���C�G��hv�qM �&ah�텈�`�#r�8�/��}�����"�=��p�t��?<�[{���,;T�kP�T�L�)ls��IBj�c.DG$�<Tt�P ;�<��ᶹbg&��9#ؕ�cn��e��N�K!���fحF��:��6�\M눩�(Wר�d߽�IB�P�$��[��Q�t�s��/��hѢ>��a^ޘ��8j₩�G@ؾ!;� r�����7�����IGP ��_Z�d���L�sn���7��M�g�w_�vas�sZ�H��ģ������Ǆ�e��T�0������E1�F�����>��!��f� 0�������#؏|�#�1�;�aV؎�f�i�P����@I�mՏ�oZ�f���;d����Z�d�2��O�	' |a(�CQ� �C8�2+�*�@LyWN��k�H`g$�5s˖�ᇿ�R�K�[�j｛�Ғ�w�[}C�
���<��������8V�=��	�h0G�Qi���cg��~O?��!��㏇�(�*k��8�YH�@(,�3;���9��	>0aGރ)�3�=��Ď�a�|���V������d�}���e�TQ������@xʁ�4s�=��Y=���}U�h(6a�ZbػR����Xe �L���0v!�;��L'�w5�Ky�)���i�Ɲ�e��1ʓ�̹q^TF+�6J�e2��K�K�����/��;�����*��E l��+��#������s^	��a�=�P��.ۭ+������ְMXH��ꐪSO���:5տN��(�kf�C�H�Z�`A o���>")�=d�X�D�M�x���;kҀ-�	�&�i!��%��q��tl
�0�����,�=��#jk߬2���.e�2߸��oVs�ԫ�?p��u���'x�Ͻ�碑.�0����~a.W�b���@��b�;��-dG*+a��=�	�� m�cUB(mm����Җ����%Y#횟}�R��Tvj���l�ޣT�Ki5���/��z��X	�V�	�9����\�{ߎ*j��)�0{�"�O��":��<�F��T�N��~5���=HF��e��B�j�G�M%͛w��>�uv�������+sZ��S��8U+cC��T��7"D-��>�����8I r�c@�;8�����N�ҹ�dġ����8���^1���3|��`@�&� �h.H!ף�z��.es�o�y���k� <f��Ec+�����!jg�}��;d=��ߪ��6��� �� �8V�^J��� ���@h�|�^P�9���w1j���"D����W��+ck\"*�#%,8�8��ؼR?����v�[�v�F�\�Z��[g��A�J�U�6&)�J' <�PeȘ�Q<c�ڀ�� a�;j}pL$���!x�}��#�-%08�Z�R_���*�ݡ���n�w�Σ�p����v���詧�뭚0� 廉��R�+��$Yc06�?~b��� + 's�'~v~,͊���7�9E�0����s�{z�?��ݗ�����	�v&&��`�����^?Tf
)'Y�;�nXA��5ƾ��|�	��LȘS?J�s���������z���a��}U�輙pl�v�\S����&8�!ܦ
۔O�&LX�� ��[�� �̜��Y`�0a�6�A8ؑTR.]��]�������f�#��
B�ٕ��>���T������i��I��5U	�4ү�����������Z�r�82A��#�	����/_JY�-Me͞�A͘�%�����|�a�ZӮ�o�SG���aB6��	c���K5 ���NlvJ��|���aV�h1?��o��0h�o��D��p{G��d�E�l�4a�9�{`��
6d�h�إ�z7	S;"��}���f_7u�Ø���ؽ}ݢ��'����F��رct�ߢ7|`��t���t�@���<w~c#ƏB� 1�%��x �f��}�C
�
��������?ݷ����4�v5���	��@�;���Oݡ�����ܻY_��{t��x�K������NtD�T��a��?t�z�����g�_Џ8�/�3���\t����xG bk�D�����t���K`0���׷���ݝ�R�-�߯3��6m�ܡy�>����/=������:h��*�K�P�.K텭���˂��5�*D�9~�m�з��H��Ox|�B�E�a�(�f��2�_�yET�\����a�r-k�f�0i���&RI�F�%[�Z���G��'��Z���~"L�8a�@���|ԡ:���	��+^�[��h��i>�����go�� 0�r��O�� $�>���"?8�"%� *@��j+�ج�.��,�RU��K��t��y�w;>�z೚z����3.V��S�ڒ�p�N3g\��SV6[��U*8�f��a(���vad�`r�~ ��ih���^Ԯt�.y�����70���Փ� ��Y}��o���U�ZJ�u�t�9����_�u�ݮ_����������?�9T�G���Nl�ٴ�����'l
��
iD*�O�_��onn�-���hB\a��m�Acv��_�4�'��wQ3��b��&,�u*~���e�ד�J]]��[o���iӦ��؄ǯ]M�Ɖ�	��a{�t�t����أ�Ӹq���p1�����?��`�&�a�AG1�s\�+k�1���3�LJYb��f�\�LV�/|�AE@�<Xo�Dz����(��on��j-_�gM�����7j���ֺu�:����z�e5�4��A�����c�)2��ׁ�6��4��]/���D_-�Woҍ�iD���F��|H����TԜy��Y�RG�f}�s���=�55�^�Ι�>$T#ĻB6]xU��}:0�ڍ>�1G=a���-���s�����:��#+�〯Am����C� ��]��%P���� s#đ�9�V>;�ӛ�Q����% <a��cʅ��ޜi�mη�yT��2U�7-��l����S8� V^�upN��f����F$k���7�G��T�{�VI��io�{1�ݖ�b�v�؄�֍��ݬ�z�N��מ��ԟV��SG{��j
�`�9+؄��\�u��N\�W�-R���"��1¶;8ݵ/���`y�H൓�� �l��zh�u�5fTJ��z�f�z�*�.��W�>���I���[u蔣�1M�1��d�^��0�
3�ܹsÜ_�j̀��������ĵ��i �d�;��8잏 ,ٿ /�؜	���L�0�g��qŕJ��9��[o�5Lx\�xb��
�d�D6�mN����1�����B�Pv�(�����xl2 0���#��@�]�B�	cv�m�qp��5�KF�6y`G��υ]<�쬑�1ݐ���_�{B���^G���:��m���s����؄{�VΜqn��H2�
�i+(��A�v�N�	�xG�D���+C���L#!j�4�Ϲ�PL�9-x�A廪7:�o�0�ՒVO��5�
��/��>��Ɩ�JSE��v��U%D-�Y�?f���p;s�p��͋`�
���?>�)��El� 7$�k��t��ǥ-}�XomD�wo���@8��>:w�܏�n�DG�ߴrQK��D�c�ʬZU�2�$[;1����!旕��sgX� \o(	Sv�84�������5RFWWO��^�u�{OOWXA�	'L;a���`�`�-w������Ru���K*�Z��6�;�*��4�PN+���sfhʔI��Q/�=�Q3�H��i*�8|��r/X�����Ȏ�F$��I�NHQY�V.	i�]my�4�u��W��oW:���fG������)��Q���Ja�V�$`�4����,X�Y�%m��k� 1��j���|M��/�7��p��zY�\�;��r��^����o��U�J���I5�;3�8�
��&Pώ����;4������ $�"na�ɞR�0��1���q�^޸B�\Y��V��W�I7h��n�}���^U�RU*KX]Uӧ�*���M���ԃ9���AB�9*����x�����H�l@y�5"��N�0�d����E��OiTSV^��t�a>aehl���T��Ln�R8�S9)ݓ��R��L�1�_ޜ��Wct��I�5�8�y�\�ak�6#�D%�b�͈��7YuXm|_��X�N�ӏ�~���+u����n�b�b�DG�Np��4�g�!W;��ǳw��ةeAqm����������?8��%������P��nP6EUa���F�Z�I�FOT�RV:���Q��;+=a4�8�@v�X�Y<�5�xa�ܯ�$���l	©���X�7*t��l����UU�Š92�w��u:餷j�}V�X�bU�$Ta�`g
"����-�y�0�dk4c��9�j��kƱ�����9��սE�|m�g۲ύ�V|=��L&��m��v�����k�*t�4Ä�ej�T�& 3e�h��r�7�c���ʎ-��8��1��Ât57/tX5SE)�YO?���=�P/���5�K���ZT�H%��Iv��sH[������PL�jmÎD��O~�`Ba��S�Qر�&(����#�m%08��li0!T�%5d�JU;���3� �f�l�0f�z�0�5�Tr|p�=sɅ����1�=c�͵ф�1H:2��ʿ�e��1q���s����L� �N��3����9�U;��M��|�'��}ͪE��0�#P'�
īIl����U��lA��@��<�=okU���!j0�r�]O=��
I��}�
9�ꛓ�wҝsd��8�����O+`LD^Yd��h�XW��f�#{��	��%˗�z�*���*aa�ʅ��Ad)�ޤ�R��@Ө�*���5%��{#h�	Ywwg�Y���f��&s	~$,�6_�q̌�ƌ>���p�&E�|��Zm>&�����;���W�)e���#���|��ի���X�A��qm���Z�N�	�(f۱m(�	W��ݪ����ڸ~�����rwO��+��P+�Q�J:ط���szm��Ʉ=` c��������Ӊ�F�v�,|�q�#��cF$0��&���p�C*vQĦS{���1Y�H��ԩ���1����G�=��W)5(��뫔X,���r98֞|2�Z�����kf��h3&i��c�5�Dc�#f��c��{̒{1m׀�k^Z�R�~�@�T5٢�/��f��+�k�c���%bVBǂ:���!(�f%�  �X�O�sN^]k5z�¾X��Ű��ŭ�m�_��U*��Jg�# <eʔ�6G�]��� Y���:f��w��,RC�p��	��e+_�׿�����7�NW^u����#�V�
Ŋƍ~��;	MjT*�$=�h<��|Ü�gBW�]'�I6>�1��6�������c��ٳA:h���0������y,���k�����Ͽ�Ug������W%pcP�����m�v� QO��X�<<v�&��M�`�<,?�-���J�.���~�(�_�\}�TNk�:w���`a    IDAT���G9�2I���ӧ' �#�����h?�7+��u
pf�%�G��q��w�z��N��A1�/�õ���0|W��Y���>�L�G.��ٙ�vN<v�����/y>���hVIs�\���y�r����FUK{hs[F�7�U(eB\=	��Y���5�xLHb�y%s=a�ۚ	�x{�qb�'� x��s�W~����&ĸ-q|�.aGG�*u��=氉'�l��|H�pt�qg��@v��$aN�p�Z�[���yW��5�2r��q�M%~o
Z˄����Ӫ���{�{���õ�����K+W�5}���jR��S�.'v9�ܙ�2irȶÑ��+MR��zW�����'C���svtt|�dlj��JaG��?�M�TiKIQ����n��ğ����{K_�)���[]��?�;�lyv5��kp�s�U�\|��������;�l���=nG�G������#�RW�f�]��[ޯ���%$cY����?��C&����N��:KeRɶ����Y��ɞn�i�1	ۙ>n��\�w��-��o�I���N�5�����keҙ�ϟ��2���5��d@�=�`K������x��44�w�"���3�p�2 �ٕ��X[��9�v����Z��Ԝ��iݚ?�sO�͟�Z��f=��Z�:�*ut7��\�t]6DI�7s��2E�
ay V@���ϔ���U]�>������|�eb�-R�L�d"ZM��[/r�N�-������F�����{0X��D�Ɇ��ҽ�1����}�xy ���緅�mӇ�a��`�����k8�$)+��|�2-Z�/��lӨ��n���{ީ*���G?����s��P�k>z��:�x��;�9�TnT]&�j%?(�������w��П�o;�I}���n���`���~o�mw_q�qSV�H�����τuk����0�R3a2� u$K$5|c;�iz���I��c�k�٫�s��wtv�Z�+N{�D�퍼l�
f��ک��\0Zw�y��9�h�^եw�~�z�-*T����<g��v�R�l0q*3�{Ad��3�-�[*��>��I�c hIo���m�3h��kGA�(�[��=F�w�~}�m �5���c���0�$S���{�!A8�pU����\m_���f�ܺ7����P18W�t�-\𠺻6ktKU���A���ܺQso����ȟ���[���iǩ��M�l&T%�M��Lp1�ZSA-�>>�d�� k?��$�^`̾��� ��cRi|�%�߻�ۮ�8a����q��Z&ӥ�M���۲WS|;�\/� ;�l��m=��' ^��p͆m��M���%��i�l,�t�N]m=����5a����懪m+W���PGw���z���^s��:[GN=J�䒌�
��w\��cOa�d�0ch���v�z:���Y�1���b��$}
��m���jp3��(ÔR���H���X�v���X�I�h�����HQ��=~{�E��ķ9H�v�r[�U���}���ѮQ�Ӻ��K5}��նi����&�ት:���u�e��ɓ�ΕU���r��j�8$��i7C���\r���;I��w�U����\�w̘Ì�EcsD6���=��s�a�6|�,�ݖc&L5@���\R��*���!�������pd�'*���+5x#(µ;#���|;WܞT�*�L����-�d˪��K�W����?Ձ�ї������?-�E�Fm�)U(:Bzr:2َ9�U��]ׅ��v�����`��̒Wt�P෽ ����''��&�W�����@̴������>��)���`~��]�Y�4i(�p,���� ��m�  �~�˖/��C]��4�Y�e�e:������������i��u�'g��#�R���i�V.���	T�2�؜8T;�s�:�#��c�F���Y&�h؄�Q�����xf0�S�{�����{�U�
�G^v�!�Z�,h��<��-a�N@8�K���[���!����aa�����l��ST&5�N� \���h�|^�öG�ap�a@!�`:�'e�舸T�A����wv���/WJ���+>r��Œ�����>���*����@u��}g���=^�<!4�`��5�9b�I�kn�[�q�$v�����@oi�P l�ؾ�a��Sj`�P�P���^����P6��Ȯ���؄��M@�H���՟\SJ)b�۽0DK�6�C�;��[����2GP[�[�\���657V4�+u�'+��~��g�������h��>v����T��Ov�	�l���0�0°�F��1�M�i͵�(f�: ��h�^��:��E0������7��7�����n�͙3��a-�~�U7�ۆ�{:�c��؄�J��l]F�[���Ïu:YU�0�Pi�0'������c����fwꩧ�z���8���/��{�e9��.�f�\��A�+�VL8SV�g��x�'�<y/u�!��˨�/k�ڂ���~�wfƣ�-�}�{���p�J=IȌm�M�!A2������w[�l���@x�I8�c���?`�j���qt�6����Ȃ��0���j�^-�m�{�/�dk��|3��(��o���n3~mӏ�@���y$�m�0����� z"��3�&�
;T,x��*���PԜ�.׌�*�+�����K��ǧ�h�����_�C4ԏR�@�U.�Sjm�1�����k�;���di�=䍲d����k��%a��l6���v�'�x��8�����${�Q�2�I?v�]s��퍦^��I�oZ�  �� �M� �����~�Lc�� �m*�6��@t��T�uvc����1w������c�=v��&�	so�f΀�%�\���U��Ù)J�M��{�Ǝ͉ݗq�Z�g�yI]x�:�R��T(R�>]o<����	�
��bZ}D��c��VL�wB�fǓ�f�m0�G0���1(hl��k~(��\�õj�G& 80VE��D�b�ۧ1���� ��18ԫv1��0��b^�z���_��ݪ�/��[.�y��b�S�,��ܢ��Ps�x
�r5��b��+µD��?�]�&��5YФ!��*8�\v҆�T�F4z��9��=�zꩾ�,��e���]
»mZ��9�y,NK�I�����3�l���z��a�"i���A�1x�#V����g��q�V/6�H���/���?�τ{�U	[ }�_[� ��N�@��1{7ͬ�w�*�jk_�Ɔ�TI
MW+9��x���o�ӓUUuJg�rw�6Y�nPkx�I�ϖW����n�֞X��)_
�℥;3)`xXM��JbL�H> �x�����g��6Ɩ��P&�>U�8��!V�X�ֲ��VD�1�}��'�%���,�Ύп��+~Nm�ĹB�կ
a�������F�]ñuu9
� �*�ej�x"��{�����I)��λ%� �O� �-�^��ܷ��\��I,ט�$~�$���t~0p��P��$���(̍�8���uu���~��}�qe�%K�����:���IS�0����j�(j���C�\����L�m�R*�jjjs��ȩ2N����\gW�g���ȁ0S�����TfK���Ȅ���P��Nv����ga'��  �`	c��M��p.�I��aA�e���q�]�L�:u�v[>��O��v̓�
��2�Q�(�?z�({�њv��Z�z�V�\h���=z�Z�^i���st�ݖ]�΃��`�l�	�bOfu��y��a~FV��7�����s�;6wl�eu���O��Z�v�Te�����ƌ�C�ֵ�R�*+5�Q=��{ϰ��{���ޤ���'O�؞h[ؾ��l)~@mY�aI:vb�J��!^�.I��e�"���8&nG�����&��+�)t�A�� �j�'wr�d`�a=\{7:L�c;�(��bU
q���`�b��$B���6�j�� Ό3#c��MS��'��"c�&�<b�N�p뢄����2�<qó`!������_�O|��8����6?,5f�-q���/*p/z�L�Ֆ
_�s��U��������=�+��6��o?�Xجa�(�D�ӄ��e���w��ή���Mx�Nz��zݞ�W&S�8��qT,�o	�����K�ro^0Q�a����wt����;� ��Ny�P"ֹ	���Ш�M ��/��!��x1��&X��6��'�%!ʢ��� ¹�G���k��'�]�`K�+0a�C���#���w���`����/���\~X `��:�4���J������}��U��a2�m��0-Pi��b���_���m��<�`Vm �-�R*t�d��*;C y]]�@����=U��/{�'gUvf�i[S6��:1�CH!�PU:�ˇ�AA �PE�E��B	5�Jo"Z�	���u�;��y�ݛ1����_���o7�3o����<�Γ\�e�!1	����Xc���J\�?���V��/�9�M�;G߳EwY)̼6�n�1�YW��ݯ�Ɯ'����8Oĉx�|l���1�
�LB��.��m
����A�o9��Ka�M-�7ӓ�GI�1aס���\���}�SW`��-"��.ס�Y]�J�	Yݫ|\��/.\ǒ�e�� $�]�u%qL�����qt��Ɉ;6@Ι����(�����g���Y�q���f�v������"�#�qEr�������ΊAXI	*r.����f���?s�!, �8�	�-�;�WX�p��o��Ƶ��Vj�7g�IsĀ�"8�����s�_~���٧���H���xI�^x��;��Q��Ր�9�9�?��!+��G�l�3*�E&f�E?��n�����OħL�p�p���[R��Ƅ���1��n�0l��x��iX0!2�\����ׁF��������:o���τe������K�������O-��|4��b��G�i�#� �͍`��)�x�|���4�2���cv��B�"K�@�A�<�aw���d�b�n��i�W(tXk���K;��%׽�Mhg��bN���9q1;���'&�	Xp�l���Ĵ���F��3y�v�r�#7Q��h����u�����x~�)����-��Il��t���p��Y�]���������M\~^��B!�O���g��j^��KznceׇRU<�����a5:�qH<����:	ܦ"�s�p�A`/vk��W��6k1o��;�2�x%A�[�S	�k������\_�by#����o!,��@R�Ϛ���	ekκ/��B�4��phqR��&K=�s��:�����&��_��5�y�d�Č]w�Ç7}VSY	���6,�B5���O�In�$���)S���^��)(�㱻ϟ8�Ǜm���e����[q���o�gќ[	�4��p5���H���^y�v5..�^����T�����e��鲛�c�=��6����(�����o��Ád9�	d�t�qqˣ�����R焍!��k����s�Q���B.��H��#W4d���>Y<G`󻓁v��0���um��i�S�Dt���a�d��N�E&78����Kf#UE�t��X
�{oQw00N)96L6K0��"�O�}3V�\�@�G)��~o9�c��e����<��F������T�0�D��ɘe��N������ۏ6�U�Ϧ❖Y��j�MQ�3�Pf���-�)�h�ùm�<�4U޳���˷��E��7�>�6T�"!�yw�&��O@��κ�g�I�):s��Yleˍ�)���E�`�M±�~�3am���ֱ���e	
�����,(ֆ\˳|�`�e��6Dm-�J�_Ѱ�b�b�$f�6LwL�i��~�3�u�Lc$�<���������_}�J�e�,�����7�4���0ٽF��׿�9�;��8��2�}Sfu��0��X�΋.��na����?����	��m[(9�{�9�s����"2!	�LI��JiBp7�JoaýѣG[�w�)�y�lxI� 566b�ԩ֝�裏ƨQ�p�W�.��ó��egJ�)?X���t��{�>�+�Φm�p��Yh��G��6cCe�![��P^�![be�N�pq�j Д�C��T�0�����C)ӈ�P(f�;{����,Í�kC $��������9b^�!$�Vf<��-����6c<C.H���]��.����\�%Ky��(����N��� eN��D�{<F�Dc�H;�sa���%���P@2�p�8S�MvW���L�������ܡQ4gn�����댚�Mn��p�?O&�+�ȟ��ʲ�9�'.ŀ�Y^?磫0��g�(_3�Y�,��ٹ2�Kõ�2�J�S�'����2i�*Y�Ry8IT"�d�o��ZfcXB,pL���'l}�Q��䇡��m��E,p#d����#95c�2�aS���8����ǒ���޸֙��O���� �,�ʉWd�>� ���_1bw\x��?�V�d�Esn#s�qm3|+|���������3?C�fe�Ձ�d�2�������"���3L�rPi^h�A�t�;�hM29�P���n�B���k�ΐF(���@g>v�<� \D<Z�[��B&�;�4f$@L��bY�$�vg���AT�[��}����t�71�yPd%0ǂ�1�x<06l�/:�� ��W�dO%�l�fs�NB1���f+e\�u;�N�عr�	XB.OO�[5�B�͓��e8qL�\+E˱�%45-� ��<i��5�g���NOfb�����j	dy�sx9&�{w&���
��W�{�F�nFZ�Ӳy�/c�9nv�n��5\:N��-��*��(9& Vŭ�T���?�.L�t:�{~����@'5e��x����:	�1B��M~_,��9G&����|5�<��:�1:ta��� �5(;�wY}���y}��f��,T"�CaB� S����'߷�%����*������q�Ɋ	��gZ��{y=�2���;v�������UЋ��t�I.�L!ي��嗝�X,�h�x��d���z�ͭ��X�.8��n�MN8s��f�V�n��9�6#�a����}�*(��wN�{��9�xѼ!���mg�曩|�4/��n��L -b~�i-�4��N8�{Ԇɐ�ߘ����tP�RϪe������3���O���մߢ9K�vʠ]r�h"�tXz�	:�r}�R������ �@eig�9&�r#��z�������O=b�$R�u�IUaIK��/�ʹl���mns s��4��A%9�ts��qV��%��>������ NĀ>=�@o��M�,Xf�6O+�w�f4�B��%�h��ȤsH�T[��6��Ǥ�Ǆ����K`�����-���X���bsk�ѷ_O��vC�݆C�*E�cP�ˆ�����ظ�D-r�<�j�1|Ӎ�e;�ܷ6�"�!�Gj0o^#>��3����������ݕv<òsѴ�(����·hk�!��6��Z{�(�l�"R��p��7��#H��fb�%��Pz0�76�p]�76�q���Yb�N�)��%����ȜĜیJ�x��У.�|��E��QJE�:�Ut��;g!>����q��O?9���4�ݳ\:��X+��ǐ);;��<�2ea�h<���� 5t�1D����&�u#�Aa�}Y̼:�H����B͗�9s(����H�د�l�N=��M]n��E����N��K~����9�x����;����"
� 2��s�>�[3�X;��ܹ���۷�>�n�b�Q;bܸ]��?^���s�	r�#�!P0v�7����Hy����,й���h��sg�Ճ�Nu�q���������>��c���ꪫ�5�嬑�T9�:��	Z4��	�?*8��꾻�d���i�jg�0S,�A"�g� g��x�5�$c�C47��F��d�+�УgZZr�b����_`��2�L ��{���N�.z��Ҵ��uJ�(|%�d�s5ҙ���V���_,���ev�5�<�$\�\1m��	^������e�����p%��    IDAT���"_�p���}p�٧b�&k"�ʡ� �L��Eʱ�b;jkz�����^�ioʹ��h<�w ;t�egS4�B���w��Ƣ���-x���n��6���@�^Q��D�Һ؜dEz�I��)�t�U���o{��L�Q��Uᢋ�ða�!�����i��"��"JQ�o'0{V+~��3��L]��^=�8��ð��۠��N>��_o�����Ǒ�U�W߄�S���O�9zc�q�ѧ���:���ɍ,�i��X���p�ݏ��߄L��G5���ß��}z�O�!�.搨�E&]v�E��T���᷿�f�Z���1c�G������kY��B9ϹYlPfr�	���^\���ٯM�M:�	´�����YSr�If�8��~{�,Ʉ�|�}�w:�h�I<���>��S�a�� Y����$#vQ�B"�|�9����v�'|����]4kR��y[�4�6�h8=����VA� �L՘i,t��yʓ*p$�e���	~���,(A�7��gJ�
���79�ػ馛:�׃�j~�Xa�:\���,Y��c��V%GÜ�T��gc��F��i�(z�^��۸&�b���j�z�q~�r*f�`A}���8��q⏾�d"�0��L	DB:G��������<Co�5��q�Uȴ-���7�o.;U�EDb$�=Ē`B�:��96���}�M�?�*,\�A�cР^��տ�F@UMK��B���%KZ,?�mB}�����y8�?�g� dM�h�?�;�\#�|����ȤCT��@1�As[�9G�~q�p��Amu�\6�r\���У��E��I�si�riԲWU)@6E����wN�E���b�^�S�������2��t���׺���6Ī��a��-8���֜4pC���y;b,��<��zd3�9]]M��B���5ho���s���}ɮ�6ဃ��ŗ�eV_U5=��҄H����$r�fD#Z�C���_q��? �gDK	��xn��r4� 
�PU� �#yh!�E�Q|2}~���a�Bnp���5�G��/\גDW ����1˰N�3�W�R�+�>�� y�G��Z%0r��QG6K�!A�~+̑�F�ʸ~�Ƈ~ءo���������=�S��;�c�Qq�a��*�-V]*���x|�ĉҭr�	�i�?�:�2B�䌎���:s��?�~�4a: x1��#;�7$�P�T�p8J���@�T��M�j���hq't!1α��\Dw8e�H?s������y1a1hm"b�_�u�)�����z�U#�m�5� ��C*�ܹ�0����޻�n=�[�a�u��̚��u���q�DZZf���cL��.�0�����O����ת�&Ç U�B6��g]�{��+°10z�!��Wg�GC�X���2M��1x���zۍЧo�m%<�ī8�UXҔC6���5{�ګ'bذ5-�z�&L�`f�^�D�
#Gm���kP,�ha��#|:�yV�����ӱ�ޛ��g�t�^|�~2˼�[l5n<��J/'�����Ȁ�m�&���r�� �x}0�0mm-Xc���醨�AP���;����X���q���a�-7B2Z�3fᓏga����Mb�m6Š����=�Y_���C��9!�R=�f��3�����BUUm�Ux���1�3����o���,"h�9g_��S���,��"|{�m���~�T��%L�����4�J	����t�:����}n�4��t��Ym�h����5�ć=���\�Ӧ���K��l3bK����|	�ޞ�SN9��f�h�p=$P��A��Hi�_g������qq�+.~%I�좋.2y��k�5ف�ε��q��g[� �F�>]I���d/2W9��Lc&�Z��������˟~b}�+�P�Z.�b�;'N�����?cH��_L�ɶo�L���܆�=�b�}��A��5.V��r�)���r @48�*��;$w$F;P��K��?C�7��.���p��Q�9?TG;��&�AO'�"�4�d�c1��d$��`.ǃ@8Z
Odp͟.�v#6A.�Ƶ�\�{�z�L�d�l�)�8�x^k >�t6�9�44-�6}-6���N��(~�Y��������-ns�o5��c��^���b�s~~��o�ek�JF��f�����ƚ���������Ghoˡ�z���18���Чa �|�e��G5hM�bР:\s��>|]�����<���hivyc����~�t:�c�>�L_�b���
??�T|��/���)�������K����V������{����������)�DX�>������Ä��_y#^}�V�y͵{c��vŉ'� I�r��8�j�Zcu=�����м�	����x�����j����Gs ��>��Gu*�|�A2Q�T<�?;2֢C�L~7�x7/\dRĺ�Ʃ���ѣ�`�b����	���=���~솸�Hā�>�<~w�x��/�0x@_��q�w�������I��o�F{:@�*�~��4�2�ѯ�f.���G<�̋h��|���Gu �Yo}����ޯ�����t�0�v��#1�n`	K^U/�}#q�V��KVvmq�Rz�߇�0�F��ɻ����DKZ�*�Đ!j<%	&������E-�Y�_�!�.C����'̰XFr1Ȁ�r�H�D���O�֌9���1��ɶ���,̇�S��2�v�c����{���a]���29� xC���!�exژ1c�ǝ�;o������3��Fq��%�s�YҒ�뮻����4Ox<�QҲ+͉;�9��K�Y��zEX�M����&g�:�z�1��`ܸ���k���������j�`޼�h�_��O9�}0�,n����%qsƤ��8��#�����s֯���o�&5������������~���/���Q��ZD#E��.~q�9�7�?.��j\����,�b��=
�����1��٧_'��$�-d���^����0|�zx������}�a1�"Wh�O�8�]c/?������tR�)E��s~�������<s�8ӢX�aqS|o~y�D��q�����?c�� V�&��[�E���e�^�{�~
�4��#�������?���C6ğ�<��ş�̉T]\�s0f�V����qٯ�-K���ޞF���<O��T~���p�yԉX8?�T�^�6�}�I8��=1�Ïq�����g��"��2��k��췿A�Ǚ?�S�>n�z��{l�_]:��/�◗�_0�)�$��x�6��.9l8�L�Ɵ�G�"5���֐�x��̂����p��+P�Ҫ`�q5=����}�݌����s0oN����lQ ԃɄ�E L��ײOθ�y��5��Ck��K/�O<a��.�đb
�$��R�rY����$1��u��� _r�wՖ �&>������z�vN�XG"�0��5q��S��7���k��7������t�Tס�.�_���k�=��:k�i���O]3���y�^Pi�t:q"����d�,ʜ ��3��w5������w_LFN0YCF�������{Ȝ<���X�I�U؂6�Jv&O�d���:�Pl��ڶ�����>���o��C�����h�^W^�'��һ����p�i��\��	S�~�s���`�� ل���;`7�g�~��r/Z��[�������x*�)S��鍨��l�� �G�� �=�������	�͘c�o��:��ʘ��t<����=�V,�U�؊ۭ�]v��By����x��O��=�z���N�ƛ����x�Ǒ�31$Rq̟7]��{wD�$}�9�v�ݦ�&SQ��iss�V���;�'����/2�Y�Яvt�>Xc�@���?pß���y�{��:}q�O�ƀ�x����g_B6�7Y��nɒ�a�15f4��<~y�o���_���Jओ����73g�#�����
�B(�h�B}�*���H$���C��ǟ2���6�}���/r�y�������OQW�a��l��y��X���6�c��������@x���8�'G0���0��� R� �@u7�F��ƌ���M�﫮�'�q9s�1���%��rK��rDe�D��EI %�u
�ZS$I���A�c+�%�����Ep$8��O��"�����~%FWP�,*��H��K�@[�K���~֡!�f�C�|�U$)�b��.���w;�?���\�H:�k�^���*K[�e��H�e0{�\�1�/e�H㵐�04�L���ed����l:?�L�p��Z���~�;�ŸH���5N3�������mI!+zМ.��K,D2JW�+&,JfN' �0Lۍ���ią�[ٌ��̌�\��<둘�a���;�Xlfu*�	'����ej.j-�!��X*ЊR��
�B�5ep�ͷڦ�H�=��[l����e�!��^��
%;�'�mv����cūo��X#Fl�q;�E]}5r�64�����X�Z8Ya�#H0�-���>�*��y�;dm~�Av_�7$��%�d,i�0�!�K�����0��|�-6Gz���~��dN��C1����JAU��Rֱ�\S�����c���a�=v��^
]]�\9�9�k�g��h�T5�z�I<��S(3Xw�5q���G]��7�7��_�A��L������,bL����%QW_�}���bNU�&)�N��u��IV�"��a��&���x���P]�n{C�1p��I�NQ�Gl���N�P�#_hCMm�eT>�̳x�o/x�i��ɣ���י�]}Wk_����(aE������H�3}G5UH���nSK4��G �c�ǣ��r��7�҄�Yeg2i��(7^j�����r�A)�H�}�9���[C�Ȅ�͙�F���ie3y$Kq˲bg��F��vێ�@tj'�%\��+Y�?�+Qb:!���ܝ�\`.vҥi���;��LX���|i���o?|�;߱z�<�@W�&���,'�o��{����|&�0M�]v�	#G���{�P���
�X���1�ic��.7�x�̥���ȣG�:��T;0M���Q���j-0v3Ӟş�x5�45�Yz�!�c�M6�D�D��ô�(�j{{K$��G�0�H�}�Nśo�D��a����hooEmM�|ȸk�YSRr������g�J��Ͼ���z޲��[-x-�r�������L�̤a�X�u�]k}�^=�C�ydŁ�ģU���N�!��1��af.d�����m�[>z�Hs~Qv1'pZ1�L���X2�x�������G�X$e���\3jj"V2'u�z��Z�03���]�[n�dCF�q�!Xk��(�]-�|ԅp�r!Xl(ɢ6��A[&�|���w��=��M7�L���8b�h�)茲�����H%��w�Y�)NX��-����kM-;��s���Zת)�26]���|�2�8~�R�E�$W�B�N}�׵�n%g���H�k��GC����s���;�k�3,�8Gi��^��p2����/>�[���c��Q*o��jy�ąQۍ��oiT��7u]� oȘF�d���E�I��aLa&x���f�>c��-�,���O3qȄ��T����yv�[�ʿWFX���06��λ����0[��w3�ъM�ooO{��2��wϾ8�cгW5r��9IYt�]��ɞdɽ�T��I����Cs���r46�d�����43��h9���&�4���g�ex����B�؆v�	;�ݫ��ێR��[X�n��W���W_�#�<jbk���q�Mb�vc�>�V�%��/:��y�����OV�&!%*��&A��2� ��;�[/&��z��������0v�]Q
�`� 7�(#,��Ӳ�-6�.���yx
�b묵6�8�H�V��4�H�<��}۞�Uch��'0g�b�1�n�e0D�����A�LCfZo�Y�ш���x�Ld`z4"hko�=�M����7��cϽ��[wT^3�>t���8w�RLRJ �i���?�g�}��	slx��#{f_�W���E�$�I�fh]�؈Պ\�s[�1���,�L�Y�$�>�E��A-�?q��@,�:��tApϹ���ne�C�?k�~?�T�ό^[�b,���ײ�gRv��0U<F ��M3Ώ�I�X�U;b%S��)b�0�$�i���IK�`� ���d�(myUO�/s|MM&��Qc��.��B����VኺS�'x�nU>x��0�d����w,�{�P�f��M��S�*���b,�l:���x5��̷B���{6�h0ق)��x3��ƺ\�6,PJ���x�W�۱�.���ݝ? ��5W��^JaWq�����w���GQ,�0x�z��P]Ͱ%��:pP��Jt^:	f�������Q��Q�C=ܬ)�"��X�,�+�t�v�w�]6�8�;�;v�
�@b��<�Fj��]�&^<��sx���a���z8p�Cѳ��B��`	",�hŜ�BM����1k�BL���z$r�Vt��/�"P���]��8u�b`R����<tޚ�������`�-G�gى,q�R�yj��t�C5)�z�	<�<#���)��V7��>h+���X�"C|8J�
  VY�hԞ�"0��S�	��Ĭ}�/�*�Q%r.�2�a�_B�y��R3!3�M2z��/��Ej��E���w1dW�fk����!���x�*�n��\Ԅ�g�6���;Ժr| �������k2'@ǈ#��.;u�׸�0k����\55�V;���>�t&�k�ջh����j���!�Rk��z�e�o�|7�)��X��s�!��Łi�g����E�$&e��5&����:�_�p \(�1v���N�:�-���5�\Y���_���NE.ߊ!��G�J]�BV�rV�c���X91~������N�Z� ��p��n�~J�r��e��E1���]�h)��v�;�0�
Њ0RD�M�D ,3EV���A{�ox��Q���zb�}@C��(�Pv ��v��Jr,�4{�|�1�.4��X����׊�S��2�T�t�rW���@ A�<x7�}w�""�b��lC+�K]�9S���u�ؼe�&"x����⋯�>z�,%s�r��^��u�g-'<׺�[��t�D�H)���"�:�i�������*0}]����~W�2Y�d¿��/~ԭrİ��f��ٓ��i2�@�@���m��紜�dҨ����	\��:�/O���f#���Xd{d����T�e�����oO8�L�%���"";ﴃ��O�r�٬�?�0�'�|��������'N:�x$R���E2�@&�C"Ve��`,w���D�=�o��g�GU���{ ��a)�"� �O�"�Z��=�-�*�?��|�D�El��6�c�q��zư�Te0�����xO<�(ҙfl��z����0�.�qԚ�������Ł�o�h֝���_�>���՚����u�ݹr�1L�4	���9'�����a���23�1�HH	B ��� %��ګx�ѧ,Ds���Ł��L� �M���+0�w�:{�,�:�6��6��G=�w?c`ٴ�$�"f�k5����x�-���{��p��6nl���	+��Jo&aD	�L�ȣTt�V9FO}��K&���bC���~��0֊�$U"\>;����h����ҤŬ�m����9߉1���o�r�y��K.���
~�g�{-�q�@�J�\� a %k�����H%hT�?`�@�Kf��KS������J��C�J�_��<Mؿ7j�����:��KC
������P��*�;�}�|���"��{��O�z,2�8k�DV�>�:چ%.>�����rf�j4)�a~Æu:)��Z�h	�@I�d�-�G{o���Uy1jv�aL�ȶ��:�߲�G]8���7^�3�<��v��z���}͂".]�[k�d�%���0=�}Ѣ���Y���F�:�k1E��[LK3"��P.IF]\��    IDATO�ܴi�%���{�յ(���61i���0.�*av���x���:���?�PTW�L
	�1�y�e.l"����3q뤛��i�1��?C�Ym-��y��PaW��Pb='�����R[U2eN�-�����:qƨc�ni���qh9�C�ԩ���^� a����X��^_���V������'>P�v�S$7?��O��O:�W8��|g�_U��Ap�������[�"+�Za��3&��c�Ǆ�@�L;�����r}g��8�J�
�����:��v$�I+9��c���ϛL���X;c�]�2	���+��և�&�5It����~�L��\CC_k�Ds�Be�.vR���R�|��b�	sF�>�N|1s�1�C:n���0z�XP���ddtƱ6��g����cx���p�[c�]wq H3Z=�:c��;�i�/��"�y�)��6a�����|wo����i�ńs�E	�w:��;&̤��o���fs��0x�Z��v́��`�\j�cA����`�;����v��Q��F�n�:�:4����x�W_S~�tu�Ї|� �ץ�%#N����Ps�����?~��{�/h�Ƞ���m���R��G�U�c�>Kf��1&v�=���!��[��-�ڼ����\��I,��4~
"�pK�>�����_�waiƄ��L�(�b�7 ���^O�����F��'�`�����U�
��b�>�乕����?��n�ދg2Dm c@��� l�˝'*w
޴
t�������BVV�~
�gU�A������u�T���d��׹x"Țcs��#)����@`�<g��aޙ��y띗��o�vۍDM�7�"�;��,یBgqmV$���v����|��6����0�5��$���='im�K$�� |{�[���f���κ�p����$A&�Yh�����:l�����&��ʭe�/F-8J� ��:�!�����|�m�PS�[l6���6p)WsN��~o;Ν�ޙf��'�����:��b���(Wi��R���@&��O>6g(+�54�[lf�4	�iv��|�"�ո���z���4�୷�FS���l�a�ӷ�1ב$�u]Fl�c�W��ioǻ��f��߃�\Á|YEp]��Ȯ�5#n����������ˌ�܃0�,"ʝ}	����}��+�o��6�Ë"�b�>�7������w���>+�\j��	&�ԭ �ى?ԫq��u��1%{���s-�����v���)Mƿ�=Q�j}^Y2~ڡ��ΤA��͔�8�?9:ƃ1�1.�"�S���5��+6�����bE}���L�B�ь�l�����v��&:�Lg�p(&-�>`�VTUV>,A�=SDUu�����QưMҊ)����k[ښ]�*5���3M\' 깱:�cîȓ
�3^����<��	�S�����0��=,�M)�oG,H!
6��Xl����խ���uD��@�E6�⅝%��*�=�v�p��+shl��64�%Y�k�i�a�."t�#y�-WQ~?�X��Y��=;�7Yk4��k�8vڣ����
�	�s9�9�)WX)� mmtF�.��"C�z���;V���Qu��#X�Y������8��J�}�O�ӷ�eY����O������ar6g+��D��Uµ�V
Fu�7����\{#G�+���+e���H��i��X��~�Y	��_���vl�C
�r^}�cuG����r�t�q�c��/��u�y��Gz���g:�4K;j��v�0����`�|�g�H	7�.j�	�e'�R���s���˭(���R��Ҟ;�
�w� P�K�"��pz�����d�K�#W��%���ʛC��7�-US�w1͝��ܚ�l�c[���p|e�	��u-]�}W1��h����z�����]!a
Q(r�3�2��QZ��}�\y߹���y�h4���	N�V&LM��a�X�av��!@��I#S]z�;k,}}�����^Y dE���Ү��U�B,��n�:�@��emB�{>�𿿬��i���X6w�������0�<�\|J���;�ry�]�.!�+3_*�ϲ�>�,Ӻ������蚻����o�g��i��@�oS}~��|�h���g�>��j|�N��RZ���τ�ͼ���:zy L�/\� �O>1_]���R�v�m���[�B�&O,�ں���\+�,|���	��]�ݲ��r2��}���X�;�騩�'��D�s��%�2��د��WW����_����9���|�>�?s��k<T���-P�wĈ�ch��y%�O�c���W�|�&|�y�حs��3o���6���4�r�����)��O o� ���=|�lK��nQ-�~�&�׽��YWLjy��
<W����8�;�oو�빗'��^�2?�u���l(��X�s�Y[%t5?���|C�,�T9����D�#T�M�$�h�?ʟG�/!�X�Y�ڴ?g���R��{�'u+3m��B�	��Z�</��k+5-$1�J�݊��R��`�;�����}C���et$��e��������|Y������q}r�U�Sy���돕�/�[lV?�?��_��+��O�8珈���	l�3�������
9��F��KN��R�,��s��I��֑�a�i%�w�7������.e�q��ޮ�F��Q�
C|����Vf��_���W�����W͕��(��sU]���"��b~0�@T���7���z��������r���խ��g�v�X��q��ܭ=�6��C�/�u{}�u��@�2�XN�P0�d`0�LqxLd��L�L�����Ϝ+M3��W5�W�����Y޽�*��e�mE��U�~oY�te����o�g�.��{�:��M�n�cޏb��STWm��L�+�%�7Wa�:)�H�2���,@ƚ�Y#|Sނ/i�|�b�H&|�E��[Ax��g�װ�Iu��m±�Ӏ���5�ʾ1/~��@i��a�(�]�|��T9〱�o�5e9pl����dG���T0^ނ�	�������u�/ouu��:��]]��t�	��*k��ݿ�wI�Xs�䎅���&��}֩a3O&�̤�^ͻxh?�B�	��|d!%f/�>_�G&P3��UӘ2�^s<��=զ�@x�E]��n�MN8s���f�R�k�jQq��V ��1�����f�a���V{�`�!��y&o�i��Q����,+Ț�
#Q;i�]u��]�۳Xw%V�g7��.��O�0������*�no�����#�F@&?;�����	�lgĵOF��cc�I��8C�&�BE�+,�E�`�`�5��B���bb�AbI<#N�K<�=U�����y ~�\�-�ܲ��<�֎��S7�;o�M=�V�PB*�B1��v�l�]w�Śpr� �U�y�BJxAܱH�Y��Ay��g��B��~rg#��L�gђ�>��w��3����*w)$�������J㑘��v�4��`����X=�� ��{��h�����@J�5u�T�u�YV�N���׋��'���'�"�Na{5Ue�3�?y�-{b� �?Or�k�q��*D��)&L�^v�i�4̟w#��D��
1�1z��ǖ�l�-�9VJY�m?|�]�D.��7�Ϋ�9�2�Ѹ�H�э�{�<�䯹�c���ؓ��m���G�?��J�p�k�M�_;uV�m�����-��.��<�1b�=����=(Y���+�4FK"'�� I�H�j����*J����ĺ�C��J��CI���5�᷑H$O>���O�V&��N:�i������0g=��F��9���z�V�a�м�	o����=�
��0�P?��7�B*d���s��hj3ou����47�ݔ�̎�,���&8���oM���P������zV���~H�Ȅ�;�<�)S���W^1��l�w4)����aGr��[}�X�/�j��v����e�[�8�7��|Q$�$�dƊ.� �A�}���� �gќ��m��Yky�]����i�ѧ���[vA*7I�+�W��5��;1ی����R5xj��A:��#�	Ҫ%L遍?�P�;�\~�pw�����3���#��� ʾ��%�p���Q�$��_�����2�
/��0t�P+JФ�K�!�v�������}=e�w(cЂg�]2r�����ly����� ܻq��#�m�b��Sb������Ǉ��?��#��7�~����y�d�܁�w�d���Ȇ))(�[�+�Ѥ'��l�i��&[%qP���Saq|�����X=��#�g���;�Зv�n�ă���o�%���('���M�GL혟q�Y�
;#vH��(W(m��S^��x6y�d�)|
�0���<��s���[/�2��Bǜi�o�/�o�Z��B	}k�X�چ<�ק�7w+^$���YQyi,�$��N�⋀��3�4�=��y;��q �w+��������d�qJ�)��|��� w���ek�gW����׎ q�k}�]v1ٓ��H���I��7#���0?O�ψ�A��Ad�����^)��O,cH-ϧ�3C�Ȉ� ��N�9A8�M�����#F,�2��%�il�!Ѷh/���N����/��q��oܕ(^��r�� i��	e��)�[�k#G�4`e0��;��q�g1}o<�!��t�I־��=w8�<�����`��Ϫߙ��Y6rU�q�qW���pHA=�@K�E�� ��{v��������"��ȓ-��s��̗���@�Cď�%&n����o�u���������ގ���b�L��s�9��
��ƃ�̽!ֲp;�`���c�=�������g��5O���]���y3r�|. �勃�}�-l� {�-����;������8h4'�B����կ~�O?��cpy����ᦩ�����.���R��Z�l�cA��ˮ30�Ė���x�ڳ�;5�/6h\�� �M���u�*��+CBW6qey��5O���^{YtgX+Ca�W���β�ӧ���B�����a�S��B+�@���
'�J��$~�	�%q��=d��AxqӒr��A4r���N�V9�q���ϻ�>�ގ!jl�2b�m��|���2>���fk����x#�q��͟8��f���r���;:2�)����8�ṣ��[����}_q��q����zt���0�l��;&��^w�H�QvSP1qW�[�r�B��Y/�Q �=%��`�)�篁/7�2�_��LE��s]o��&8ꨣ��&����QF�����]E��u�]�鐣����'Ű5ʜ���v��9AX	�Hi}�w&�͙7���,����Ϛx�O�n9���5�1קq&�5F�!��n��6�g���ן3&LM�J\�㖄A@U��&�@���]L@��ɠiV�'��� ��F�X`f�q0��@�m~���|2a�t�	�Ond�����pvt�X��B�t�DZ����Q	�r6̐����	��-���?wk�OY���������Ĉu�w�u@�r���&h0B���O�x�	�%��\�#\�N^-iʝq%�������!���Cak������9G����.�J�XL�x�ğvktkG�Y<떪�f���^d���18`L��m|:�S�J�1a^w��yy��&rGVlވ#�D�A����$�g��[o�մ���ƍC�^����<�b�<��/1�Ck3S.��q�h�%O��w��d�aW{�͌��	I���6���������_�{)�m97�^^%D}�+�j�U��/���c�=f�!��W�ċ�������R�$�aZ��I	hI iE�	����+�1;�x%�q��M�L���#A>�����v���3�l�s[�y�H��Hk��#�8����7_7&LV��߿Gș�U��w��F
B	��9m�4�9�q?��Qf޸^*�̸=?/��/��$`70}�~�{�i�1���v�i��[	�l]����>i�)�ɰ��Z����uG�g���(�9��Z]�]׷,�^�����ծ���8��LΤ5L��+��{�a�7-d:��������ә���/j�T�A�O�ϑ�1�B �02kFy1e�5��q-D���	�׽!j������ϟs{u{�1a֎�]��~�j����!Ӟ5�w,�0���
j�@J���\m$�=�`�.F���Xڎ��aFI��/A��#$�|P4T�G�+��Z2�=�uK��O������d3���b۩W�2;���_�u��d�����XU#  ����-"K˻>��I ��</�</#�ԉG;��~(�Y��zU�	�0�	Ԏ������<.�%��\"p$yLS�̡R��5�>f��~��b����h$:y���u+fg�>?�T�K�
#a� ��$��;`�m7Ō/>�������f7B�T��2R��<�
��	�a��<yS�y��J���Ȧ�"?�~�̕��#��PcE��j�	���;`e�x���.�l9��٥^�Ć	��Bgw[�-Hf;�կ�#�*G@ �*������Yl�Iv�'d�
����U��N�{�)��}衇h�5~v�t\�W>(���+�e��~��_��&��A\2"���0U�̚�wx<5%�����ǟڭ �s��̺���UB1(��1d�:�k�=PSW������wA`���0��@%�̙!&|��ݎ@;v�X{���u��-z��yY;����2�H�2 ��բ��Z�.�
��9C��|��~�����׊��� ������,���_u~����X�3���yN����ԕ5�c+ոJY��{t�}��Cɒk��	����,"�u^�{&`�ES��ڣ�I����}���x#���)�-w9���\�`�*�^������U�x,�(�B��[�w�}�8o�O��n��!�F�q x�����(Cpp1AmE�9��E��jIȾ��:Қy��c����K.����_<_��@��&P��(˲��(r�J����VԤ�(�ӈ���C	���x4�I��A��kH�CD�Id���X�C�E#�J:3&�/Z�q%��Ǘ�Rc���{��eW^����9D��k���/���l�%���&&?�0C5S��<�N^�B�����ɱ�qP'��b9u�<����9�8Q-:9p�hx,��j���gxG��+IH�m�13gy�^����]�@�/E�_�-eUE"-���|1`ݏ����4oI~�,�"Q�X{�n�߅ߣ��`��c^����sI����4?Ck����� ����Ngc��M�_� N)��=�e	0���%��!G�|S�6�(,Z����<_�a4�<aw;f���|fT�����r�G.�E�=��C1f���drvQ�UGXT "vJ�7Á�.� k�&����R����m�8��=�<���ѣ�L�����"�'k�æ�,(;�J�!�L �s΋du�]{-$�r�6��@��A�G��C,��T, f�='i�a�)`$�L�5(�R#	�"q���b��/���D��q:�GhN;&�tj�9?R�c(p)?���
,����n1��k% ��Zl��$�Ȝ��;H��.�w8�A_תI,�����ܼ_��.��k��<�ǿk����Y�k3X����k�����>��L�x�zx\���������� �����5�s���9�
�d4��|�o���ᤵ�Gh�&'`�>�(mꚣ���_�y:�&L�`>'1k��X��n˪#(��h��}2
�X���#��$�3=�_�Q�xn���11L��1�U�Ԅ�Q�gFK�H�!��fQ��QU�¨�Fc�-���4�$-B�!x��#L &�gf�2�v7�؊���:������.�IC�&�r����	;.�'�MdO����ۻ���^�߷J�,b����kò    IDATA1ӌ�TD,( d+ˠ+ҝ�n4@�!ϱ���g�%̚=O=���'J�gsK'y��X�A���;ݓ��d>;Hs��4bv>��ܠ��yl?Xݟ�Z�:������E�+pҵ�!�ϼ䑖�������siQ�㦅�MC��B �3>ȋ��z�U��[<��z)�Ō���i�����|K���;����9 ������_�;Z�*1@B��?��dA�ei�iMi���~�ZW=?րa8�ψ��+c��\</}G��~�9�YqQo�~�$LY���y�_���)�L���\�VF]�4ymd��+�?��12��f mR�#�s	�t+6�܂�'�ȧG!Z�DJQD����@8Dd�Æmj^Fޤ���<��� ��:�-(�s�%V8�v]NID&e���������gQO��gpZ�2y,d�l/�#UUg�m���5����>j�QD�,b�,g}�|�bD�A�|�-GȀɎ��A1���$�u��{к�*J1̞3�b�h��	�st��\�߹�k���$WcC�6mP81C�r��g��r��4�Z�3��bx��Km��p�	$C��\2�x�ƼV�u���d���g��|����Q�h:�3c]��bi���,&6-0��ߠ���%	F�6�y]<�����1jc�t��_�9I����6$_,_l�1�$22�Y�׿�u�s����Z/��R3�5F���/�[QQ�L�o�]�$���J\�u1����\���c�g���f˵ 4��q�2(1�:9	²��L9&�I��aj�G���ɖA�-�)Gt?�_���5����H��cH����e��0o�L��7����M0	�d�d�
�֮�3�b�.ԎD;���Ŕ�(��w��9��N��"�Cј�-���nM*���$�!baI�?A�u!�p�B>�agA���l4�d}��]��a�D�%��ېˤQW宭-�-gй<<�G���z������)U\��@W�T~���h�*�G�\�W�'�z�o ǌ��.m¾i��A�����'  �3bt�~��Ѧ�"ޛ������R���6+͛J�Gs��)�S�S����޵�h��f�w	��}�XkbYSX?#�Q&�/���;ǘ����܌8b̫��y�U�r�9
@}k��'�+
��:#���ճ��7�a��w�'��K����l��*�Z��z�x�}�!�����ƨʣ�<���K��DC��嚟�&�{Ձ��ųn�J7���g=�"3�J(9�9k�IMX )-�T^��L�@@9�r����Ap�5(��q��C���~�>''���ٺ�I�'"�DY�ǙjټC2ՓN8���,�����y�GrHF��GX�����&E�"U���G��C�A� ���g�m�H.��]{%��i)p�8�b��G1+���.����)9F�?�	j��y�1�D@����5���O�_ % �=��@Z�����{�b��"y�b�bx�C� 4|KJ��a���MJL�x�t�bX:���Jc�U:�ym�E)psSVKG(�')H�բ׳�����32�}��e��� L f��ƘL�a��/��Ȣb� �0?�Dd�g��dº����>����R!�3�j���H����Ot����";ڀ�1K=W�O@��#1�H$r�����n�#�ַq��5��ѥHj�t��sH��h-��J(�d:�db)(wPj��G@�7?5Ȋ��3M��	[��	�<f< _�^:��qmU
'��X���!(��D��>F���R�H�@8w����W�"����*����ǀ����&j0{N����6c�,���uf�UN����1����K���D��4`91�zeJ�C�����O�e-Mx��򀋭qb��3�$h�Y�(�c�͚�D��1�{qI���6�JYC�$�3�g�'SK����(V� �����3�ߡ�Y�RR�\��`l��DF�y/=R�K�b��d����\��~�z˓���x�rF�=锲$%}h}�F7?K}���63�a(�֒,��7�	��#AX�Cf}#2e�u@X���!ه��¼VE�p�@+�����z��X5�-��{�UVI�M��'vo�9�	�
s�)=���9�	�YR[��<a������;b�S�����0�]�L����vP���|M�Mz��vYǜ]�xf���֣�͵����5�Oŀ|R���E�0�m��wA��;s:��F�(
�8r�v �}dP$k���9���;��ڌ�:gfs4��"�ܽ���J(Q�F�C�z��ۏ�������q�@I��u�x�g3>�3}K7�Gm
��٬ed��0rYT���1����v0�e1b�9��tJ���'k����u7���6b���X4[� ���,�5p1hް+�*IKڈb�� t����dN�\�!��y)j@�7��	�f.V�{�Kf�Sg	�Z�҅+Mf�:5S��� ���6TW��*�z��n$6��9�Pda�Mv&���̈� O<��������W����xɊd�e"�2���j`�0&k��W]uUG%2����,��{d��X����ؖ,bޓ�
��0a~VdClT2�oai�hu�)ʗ/���z�Y�֗|�o>i�����]���~���lp�E3o�˷�	3�@XrS����v�x����Â�l3q�0���C]*@�Ў�X4�S�ZQQhkrR�̲� -�56����꾨oX�d҅ �-�-�݄L��h2���3�dA,�W۸HG_A���=)sđ�߷�*W_m)�A����j������'�����Ҏ���(����!�T}�r�T���͆�[v��MNV�z!� N�H��1c�
{~I�P1�
�z�.�b���A'3W��En<b6��8�`Դ�V���E2�� ɾ�D-�gs��|-�s��&��Z�~��YM�m,0Es��O�\9En�ǝD�����;��$�Bi���"�K a>�L��=��ö��6�(#q��Ŧ۳�Ɯ��ᕱ�}�	���4$x�R>[�6
E#�|�w�H�R�u=̲*�3j4��a��>�|�$��lvQ���0:�@�M�ϔ��b�e͊l�֌��"l�IW��V��/�7�,DD�'��}���ϜT�k�b¥0�D�A�(��A��e3EuU-�%uУ�?���H�J��H�rX4�sZQ�(��m�D�\!�=��C�G��ꋆ�� ��H�c��p!n��f��-b�bQ���؋ǋa��ߣ5)d�Z�7Q�z8����t�*M�|�Y1`�Ǥ>�|n}�,nnǀ�^hY��h�X�HU��WU,�����"[4�|��OF��� �����R\�t��i��1�`�c~�,�)�2�|�B�&�P�! H_��%'��㎎��iI ���L�U�L��uP�%8��әK��7�LXlI�?+�t��zv\�L���f]Ǟ�B��g��ڷ�$���<�A	u����l��{��A���� ��mDt�K�|#� S~��6��$KE�	�L��%]��Ra������ޞAX�`�6�bǝw����0;X�`��'�F*)�Q�����t�k���. WFW�� ���u����n-eI&�k����r���'�0�Z�ԆY������^=q�1G����@8^hÒ��5�G2Z@�o��٣c/��(��#F��xOdKI|1n�<	-�f$���������K�!�Q �Hզ��V�������=� �4�d�z��"U��d�C��G>����q�K/�1S@CMo,X� A,�h2@��|ɠ��ȡ�6)Wys����Y��-�J"��$)�D$h�*١X�LaE H�g�"��Tr��tlNx�:�E�����@�lS�"8x���#��1|���^���f>ٰ6 9}V �}�Ii�78I�E	Ѻa�[o�m�#uM%�܎��JX�F��f�=0hض(ī�s��{��A�A8D*��Ի��{o���C�TD!�6&�.R����PʛdUcq	�	l�Ŗ5f4���s����'v��|�F1V�JS��,	��P�Ed,O^&\	�����lwY��}"�췒i/���~��ğ��8wR�c���4&L.�6�:���%�ƀ~8��г�B�b+Z�A�e!⥬1������0̣�h,�S
jM�F�~��C.Z�s�b򔻱�y1��q��gMPR`̲ix�� D)(!oi��tc��>m9$��PM�:,!��S���P�GQ����x�g硵��d=7��\�R�����L{�@cƬO0�� �"$�e�E�i�I��h��?���xb�2��td�<.����c�]���`0=�%���RkQ��x겼F��S��xV�"�&`�$XW:_�=�`��tA����w�I7"t�^�9bz��kT%Sv��=�gϺ�&YK��JƐ�ŰU����2��8���=_���{�m�Y�m?3���G�rS�q�ؒ-۸C�B	�I @�!���mll�d�@(!(�dzI���EN�Ќn�V���g�������[�7�JG���^K:��=3{�-�{?�S�(�jT���$Km0j��;�i���[�����)�T�6��[��p�H��Y�Ѧ�����g�b]r���P4^i��h)��D��d��[�uB�u���2�� ��2��Xnx�b@��k�yӲFG������i�*�:�vڭ�W��s֟e�}=[�	��Qk�LYbL��U�ȲV�*�)���s��Q�������f^�<�ݣcv۷o�Fc�z��g��LN9[ъ�J#�f�Yg���bv�،��Wm�=�b�i���k[�8�Vֲ�8��Z���������3h�S-�F����6�w����A��G[Pl	�n#�G@��U�d�3'�z@C��rm9�4��A?�Ctar#t����hRć�#�ع&Z,q�8��Jb`�S ��B�)E:�9F;8������(L�}Ӗ�V��`'���g�� ?0�,0a��jZ��n3I���m�IgYr��7�1��-+l��JT5k�����'-{�v���oي<�z�9�U䈢�*�~@�RK: \���䣟d���lk6ˆ�d'���|���W�򕞶���G:0񼴷�a�ݖY7��!_Ch�u����1Wh���/��l��B�|0WB���8�p�Y��n��5�-�Yy�~kc�Y�6�Y���L��t�1*'�3Nw]V,��-'\Ӱ�����3]��ZM�R��d �d�֎�Z1!�����۱3��܊�=�vD�� Hcڦ�Bt�U��HR��+�?{�:�o����,�;8;�-b{ۭ���N���;�� D��Г,Sق(�Pk`
���h���*�H:3��}J(@b ��������
`ܔ+�a���(��)����a�Jq3���M�B�V�ݚ0���=�^��ㅯ!�o�z!=7��g���C�����$ɭ�6����R�X}��x��O:�F+��N��.�D@Q�(m[�N�l¢��nw~�VYfլe��3a䈘�R���zo�j��ѶV#��Zݝ�ĭ���XgUl�pᢧ�(����i;���B�*ڡpt�cN�7[�/6��~.�\���^���΄	Q[�}��_d���*hmIl��?�f�Ǌ��Da�y�H�(v�H�R-�E�7��DY�'����L�u3��jQ�|��#�05<|$|�����XEX��]vb��Y�=y來��l7��6�YEC�]S�Z���^9l��%vOOb�굶s|����h6�T��λ��{���#�p<@IX ��*��2ay�(̯�7��	��pi�������*��sТU�[�\�ܫ��Z(X8�)�DV2!ll�%�P����c�=�x�M�h+ŢsM�?2Lx� $wռ����m�1e�(�f޲��^Kk6�w����*ǜbc�A�`���|D����ylڶ�ل%?�7���;�*ʭ�6�ؔ�@��U�"�u��Z�8��k7���h�V�pPJ꡽�H>�l�E�Z�X��������ąLx6P�n���ƈ�,#c�s��m�4�r&�_��w&��*M�1�8H �JR-k����{�e��A���L���DE��Jkd�W ���L�[9[掙��s^l$
S�xm�E=l��;)��I#��rb��Yê��f&XےV��%�Ț�������M�׬���S^��E�Iu0�T���������1v����Ģ>�X&�H)��b�ۉj"t�AP;���0����~Z�q �$�0^U��>�~Ђq��P�ó�F�@E�1E^���LZ (|�@ AX��3�p��IN`�y�驤XSN�p(�~�?�Y~���
�iN�L�p�n���F���;��;�b@8�f�j�[W�9�@)��M;,����̏�k+Y��/�ʢ(6v�a�FMw�E�;D K��$�Z��l,����Z	�G8�e���(Е�p  <���3�X�@k܆��{A*A���|�;ߴ~���K����}��lot�����=zzk�6C�Ll��aI5�v���bbk2���H0A�x�Ҥ�t:�I���8K����7e 1��/ ��F��bma,�B�Q�g����N�%xiB�Q������#�2��ʽ����,.7 �m�V���p��y .�//�<�xFb�7���qd�8��$���#v�Lj�b����641i�ֲUa�7�'�nq���m]�Ҿ>��ݽUk�$����ε������w�i���@'��{r	��")�[��_K�l�?l��
�(YCq���tb")���&�⌹&�Z��(B_J�XA�@k��8�c��rM ��"3���9' V�c�.����yV:9��]�Ŝ��z��"���r��s: <>1j	�0��hV�]�j;��-;���[#!�0r���"����#�~�&���3ូe��I�Va������=:ك�� B�<=ȭ���hi�b�J��M�҂$�J'�g���CR\C����!g>�J��`J�	�G����u�	VI�48�8�q�g����3g$_��$�ʢ(���W_��e��󪧮ڽsc}rt�(;k��d�U��i���� �9kPiL�T��=��T:���PcQ��������I�p���|抛�(�,Ei�����\��+C�<.0-�u0�D^����ck�2S	05�`_��L,C;�K������+>i�+^]�ZϮ���ɦ������)[1=i})Y�5K���"P뵑�j[�ٿ��vgod��56�hYk
�m���A��������1��O��b�J &}�s���9C_P�A@XrD��uX'ז<!ǜ��ø���}#9���o��J�a�B
��@Mǜ����M9���&�x��yf��*�IG�� |��g��������y��Ƭ�vTV�aϾ��Gg�!�b�UXЋ�9���r��|��;�a�w�����YA�R��m�3_�԰�,C+d��� S��?~�l�+Q�#�t�<�,|���|�����2q 2.�����bb���"s�EZ a�2<��5TIN�͵��+�w��qM�cT�L� PO�37�|�O>��=Ky�y������ؽe㊬qN��0vֈ��5��&�њ���!;�<`g�X7!���r?���`N��w�k���^��luM]O�Nb;4��ϺW�����S������ߙ�Ej(N�"5����e��bLg��'~��LlX	&3�h�L-A���Ľ�!Qɬe6\1��kϜl؉��Sǧluc��r���qݲ4�
��R����=X��=�5KW���f��F�z*U��11:fqT�;����n�>icͻ԰e�#0py���{��/�jCK��`<�s��ń2�=d�jG}�~���u
�	b� �r�s�	k�Q<2 ��&��Zs�ZLx)Z�Ϊ眹��䞞>K�G4��k��7�m�ն��Z�l�>h≉� B�*x[Lzs�ik�qK������_�a�+B    IDAT:ά�Lx���.�
��y�c�ѕ�(�q���\"�]�2���L�tiG�!]Gc8�e����g��RҖ�<�'��3���G��0Bf#�r��ƪ+�xU�6,��kHW"��-�c� ��`�9�.Ϫ�'�_Z��o-+��Ʒ<}�ևoYg�4[3��*mt��ƛ�6�r�w�8��}��	D�p��aC�J(�W�dV0������En>��shl�I��ƕ'�c�NM8�����:&�âZ���2��yf5�s-�w�Ee�����8�/@�-k��������<�j�bY��n6�Iw@�՛X�J��C1j�6�vB���	[9M_��Yw�fy�I�j���j�eՐ}�?���m�g��pD��(���^�!;K#��]w�=�����!��Ć���;��X`X�'lsZ:�"#�%-�0�r����s/��:�/9��o�y��&�D�$��!˓#�+:Bm��<����WY:�p�U+�r�M�ŝ��l��$���yVԥ��=QݶWW��g�o���6�5��}�0�p��r&����6v׷mMlVO�	�V�p��I�ZRK<��,I��9B�/fZ��j8�$H,�I����T���F�2��!��31z��1NȘ�KV�|f,���
��(8¸;t,Ϣ�x��1a�; ��8�.�A���1w�7��ۧ�z��B�~>/�Wmߺq�=s6�%Ӫ)�vf���ο�v��s<�3�"N:_� �י�Hc0�y��MHb8:^�N ��_�r_� 0�I�ɤB��%��ΗY�Ux�FaPc��i� �@z��ib|��ꕒ�Y��u ` 0�zp��9���{ՙ�0/t0IRL!�D=P���P�E�q�Z�e���(�ά��6����q��N�b;zt�V����ܹ7��"u��V�j#q����G��p����nzl)1�+�\~ ����羻|��.3�A�5�e�p�$=�A�R&�,�V�VR���h�0i~�@!�HÄ�@Ӷ���9�c! sK�~�P�8TB	Yk��X�@DdA�SCLXKOq�L`b��)��n�f�Ln����B�Z�z�e͆ō�����ڨUmGm��~�y�>�D��;�x����<ށZH������6qwᘫ�g<:u)��@f#���d��#3>oD���n���]�նZ��8u��\%iHㆶ
��5O��c��}�o_��/~���\���}�+_��~����N�*���T����¤.R�T$���*�B�,�|��jn�xd���7�p��.+?��o�ڑG6V���'���i�0L��S��_~�m|t���>/����>���19�ƈ��Y��>`U�+�6(c/zы�)��G��e�]�E]�������*3J%�h4�<��I^�:#�2׿�,*?�9l�� ���֜�4K�V�&�jN�X��
Ḻϕ܁עj'�|�#�^�Ɏ�[���n�z�)�@A�Z�;J(��<@��8��Jl��{�Ln��96i�hR|���fI'�8��Zݶ��m�����F��A�k�SO_�;����B���N�Lfm��b���e *���{���߀%�(*|M�H *G�E�����9��9��7,,-Қ�_�V&�駟�u�x|�,&l��(�M ��ϸw@�	��Z���!'�8�:���d��C�Y�6rWR$k G��i�*��k5��-����xT��a[s�k��X��P��RƓWHB��2[�OYv���]�)@8���̤3�F;wn7��q*�t�Z�f��Z�W�#���!�VO[sjW����_���ojk��f����ox�k� -5G Vj���L����m޼�ﻛ ҟl��6i�3@��f�ݒ��?�	x^���Y�X�p�e��n��e�5����[��
��v�QG���?r���w��o-��{;,��W?5�UޏI�C���(���(]��X�^���yN;�E4>�b&�����B���U0�7�Zq�p�6B�2�bxp��^�[�j��֌բ�Fwo�tf�z��5S�	(N��׏�#��_�j�U{V�>s�nY\�ѱ	V�zO�)�ӍbK���8d�,��
�+�<ڵ۞2cvR�׎�lZ}|�b�����H4-gq���ց��f2������Bz{|_;j�o������% ���X��i����l8F82���Ԏ��+��\e�J_�0�BU��b.���{ca��6kr��z�#��Jh�,�b9>a���l �ǜ�qó;#$��i�B�pʚyX�ӟq��F�аM�O�Ӭ(�Z�I�؞dȎ:�\��z�M��m
*��E�G�,JS�6m�w�n{��^'� \DG����r멱04,�&V���i��}���<��x6��H��L��]N�l�7~�7|�-��E�J@ZEj�[,��_z�.�^1�A�w�ĩ�'`c��������Y0CkJV��Kƍ�+�2�@̳R���"�Jy�EѦ���=oYv^���[VX�l�S��s�s�=�%��w��_���Y���		�0��L+���xp@g
��AC2�1���a�����}��C��9��h����Š��`>��a�l�]z��G���/�'���&���q�͌�X_5���������C�En��cK�VZ�w��9�ҨϲJ�mٺ��vl��`ș�4�d� �}a@ވ�	��;fϬ���k���������ӹ��"���Jl�(��������^m;v�q�kR;��f�w//L�'֣	"�U�}'���[d�hb��É&&$`���'��	�д-�v�0�K��5fd��J�P�eq]�h!���a|1>���&���Ҹ!I�()|d^����p�96^�hj�8��{��W�cםg���)���L�2�"�-�2�[v�7��v��CF�JɄ��[����'���S�̼��I��r���g{�lUʣ�� J �:�SI��A������O(,���bA�ve�/��kQ`�,���2!�n�G�w��#����y�+�����uñ/i�-��<��[n�ſ;��Zqo��޺� �&�r�#W歳(̀���+m`u�}�;���W��a��d����Lh|4���Я�6��)��P��.�*�'�U��?�4���ц��|zp̙��:�T�V%޹�Y++6���^i�}��OY_���b���ZV#<��"��`E�,i�YT�V�g���6t�S�	�}�m�۴i�kp}�U?�A�>��ĥ�I8{ r#ʭ��cy�i�Ql�񫯲��,I3�խ�h�C��FaS��Ib?ٺ�>�7_�Q�SkuOÆ�T������r�䢋��O����ov�e�+>@S&?�$&JOz˖�v�Z5!�N�<���Pp=��U_jr�R�0��~ ���|.0��%	�����31D{hR
�%o�����H��zv�AD�_��0{�|��S�*���l�ն.��N9�,�)� �@�"k٪,��އ�����o��ﱆR�0�"�O��S�b�؉	vN<�?��Y������7�f.���~�ɳ�|��ޞ�J�ô/ɋ7ݏ@=��5��7J�^y�΀a���W� _|����Ӯ3|���4��}��?A�+-6�2��"b9���X�`��?g�@�Y�J*�[n|���� L��ac[7�&F�A�t�;�^��+m��#��;~�����(:����3(L7U�X��ѐ8�ІE�FD�{��^��0� ����]t�ׇ����+71�@b&ZqC����o�Z'�b���H���׾�56�_��9a�q�vo�w[o԰zJ�Vj-*�Q!")UL�v\���[uh��}�5}��^{x�N���M���E,1��AQ��zl�G��qbc���]��W�ꕫ��V�p_m�\�E�-����s���s_��MLO���a��ٕ!q�6��"��9���?�R�ir1�Y@5�Hb�$��N���`�i	`��@��� �P؟�����LL@���/�R��f�x���*$�iBr�7�����P�ǽh�`�`�!��E@4S�5�,��Tg�����}bi��.���l��ô�
Ql��X�S�ǿ������bl�n���.��-X|faYF\w!�M8&^�s�C��������r) �͸a�9�?2�{ �ō>`<�7�^��=��p���M>%�@�s�0�9xE8.��x�,li!4�j喛��ۖ�׌nEv&c�Y�<�^���m߻�v�O��-�='��	;
C�ԑ|���ʢ�����'?�4�������C����װ㗼�%�z�������WZ�
�I� �k_w���,jOZ_Դ�[���3�,oY���WN����.�78�i֎�����m㭛mz.kΖ �a�Ԟ-ct�I�{ѡQ��e/��׮-*��5o�^ �ÌjUkf�=�Ӈ���w�w|�������0��OHL@&b�F���߀_ ,p-ڭH�`p�4%��Ľ�ó^��	�Ra.��0����ώ]+�HzF]G��k3I s�0�j�r4�Pa�R�`�O���-a#���cR}�A�>i�ܷ&9@����������j��6�(,��Ͽ��F��`X����	5qa*;[����}�KvםŶS|�K!!x��$��\ �yC�Qʲ[�AX}�O1ae>���L�s���H�ā�ik�,������Ɲ�7c#S�`���i�a<�	��5|�w3oX�q�M�ZZ�$���׽{y�0s�[޴*J�z�}v�ΰ�/��~t������Z��0/V,4��ix
@�B+6�0 h:�������h<4�0e�yp&:�R�Ť�o
KÀ<ڠ�-��R��e��j'�NF;0�g���W��@ݬ1a}����齖M���j��r�mO)�=��Mm�aFT��/v[>�ֈ������#�3�.G(O$�lM����	�31�/8�<[�r�O�Z\+��)Mo�x5Ҷm۹�n���695U��E������	�~'�|��4O7(3��7���a��'&$읶���/Vǳq-�$\[{d�v����=�هLD�Tߊ� ��������sM�	��XV���Ua���!2�CV��@ L��D���}�z�^CB �~�m�u*���*#�������I�:ŭ
^$���ʨ�<���۾ioy���2�C�`6f�O1aL�n�%��d.�{@��B9��º�����M>!��,�ZHO�Ї܊�8=;�#9��4Db��z����g�a�ϸg�k����/
�ݺ}���fd��w����6,_��#�<�ЦU�n�iLu@��+.�0��V`1at~W�Q8x�O|��	 k�Ya	�E`R���/v�ba1���\@��]8K�9�8����u���V�,jLXo���	WҦ�F�+��<59��F��_���Ҹ�ޱ�6}�3%Sͪ��@��͂	�l���SE�U+�}�+
Lګ�� �9,j�T
5���ωC�V�l=�pk��*q��Ԏ\SN�d����3�8Ma�:`T&c��,_z):.\��59��2F�L��Ư��1�c���Ɛ@T��1S����!��$�;iC�_1M}�x�Ox_YWb��a|b��O	-D��g��j��	Ÿ2&t�.��-��νV��-C�_	w[V�H���ń�����aڌ���:Y�a�� �d\ >K�v�%k��
4��|�!t|���j/@�fQ�V|/�@���c�nYv>��p�ѣ�l���l ��pʱ'��_�2�#��.�?ǔ�I��!�#@�ae�sF�&���ԧ>�lW&.ǱZ��ot�x��������W���>A?򑏸�,P�х �s9�y��)X�<4�o�{�ڪ�ׄ{��3a4as��Äٷ���គ�c.��n����mőO��#;v��[?�ż)��p�	�Lt��� �Yy�Y�t~�@���s\j�r^4�g\s�]p�|�l9�rϚ�j��ݤ���`j�#�qM�E}*kF�mh���� �q�Z�E
�C���|��o�/���5���u���$����p����I�P��2?�ǋ���g�M]HZ�
��X�0�Xp��pұ�R"U��+3]V���@x�L�@@X}���0a����|��@D% �<#�'�g8�y�(EhgA�|<�5\�4� 9c69B�E�!�q��!�@(G�yފ���_w�ۗU����wl����+��1k�d�yͫ��[�{?�ow̱Zs�au�&��V"����F 5zaj����@f%�-˩�b���qڠ��Z�tP>+�+��a��q���Wmh��)뭴lǖ�,)@��o�ʆ�"��� 4r� �n=��Ӭ���D�u��u�glz� 5��o8��{ͤSYɒ��{�ܑ操h�>~�E���K'���U��W�(4dXb���sorӳ0����Ҁ;�rɆ�������^}�1��NOw�:�Ȕ���p�$	z-�2C��!h3f����P:�:z6@͙f�8$���P���"8� ѢP��]G���i�Lu"��!)��j�7�T���(U4bҘ���q�X��E;������4a->r��Mń���&y?�#�����4a-���M=����N�ue�9�܀#֢ȹC�~%>WʱH
 ��S�� i���p� �D��=�E�d�j�z˲���+޲y���%D��=C��W��z�k�����5�a�@�ۈF��Qd:��P��TMڏwS��u�Nۮ5��q<l�kʘ�M@ŵ�4[r��pֲ��~{��^cCu���V�R�������Z-J���A#1�%�=�Ȟ�,�)�^���a�ꈧZ�j�Zݶ���L� �g�h�ζJ��:@�v"�j[S��平&K�X�5Q	.c��}�q1MڃDwv� �C"C;�m!���dR��@N]�),g��_��~
� B�T��7�K'��hu�"#6%G��s����X��� 8�F�PH�>K��؇7��ߴ�X��D@���;�̘�Á^�<"����zO����e5�m	������3��� X�c.4�Ŧ�A����|�#ǜ@X�,
]{� ��[__gh�n�ǰ/%)��V������lN.�u����P��~�2qÅ����>��4M�7�x�[���O���C�����t 4�f�yϻ�.�������'k���e�,/nN�U7@� 4���̀&��<MT~�L���|Ql�L��W���Nȑ:[����V���?蓂���<�.��|{�S��;ئ�I�ڻ�c7L�R�<|�)\���Fq͒Z�E�~[uؓ��/{��s��w�u��~�h��v�ffx�a@T��$|��#T�M �-)����ZB�u2���\���y�P:'dܳ�е:��s��_��^/��K�!����Z����Y��X�B��sHz��bބ㑬:K�`�ra^J:�3@�^�x�����U�_h�.�M
g�B$��H�S"��o@����c �*�\��9�ƊC�6`�UeG�\IE�0E���A��_�Ӑߡ,�馛n�j�Ax�O7�Ό#GD��TQ;��g�%�t��{����;;���sS�):A+4��F6��j�@k�db<�[���T��*���H����>����B ��Ť݉�ʊ]*�w<I����nN[N	 1kY�R8S�{.�+�����Ψ��Z;K�V�əF�h�P����1E=� �uO�0���J�G.y���o���ŒP�����<��7N��~ ��|-|�\�o#��ZES.����4�	���_$:��%�%q��x���g�TVQ!��3��z��\t�ԅ�d_�H��/D551}q�N��L1S�E�EDa��3�2)e=��+W�k�cX�<#�O.T֕�E�7�����e-�^�w�����s��{�����U����֝b�^~�mߺ����d�bt;*$�����y���`�$|�< �)�H���f(z��>�1�
�g�h5J�����&���)_���l�AW~�`    IDAT�d����j������JU����b��)Oi��B�����1�Ez�I͊�d�N4ݟ����췀S����r~��&�;�ׇ��������Z~��@�쁞?_�?>+,����H����^���C e�IǗ�S@�q�����G��F-0���_j�b��f�V� �A��3��y�	��_��_v���)A�$~!�D��z�~$e*� قci^�K8���H!�'B��k���S�_�� ·�����ea��_�{��3��R� M8����	§�r����}���ǃ�)�W�It,l��A��8�b`��e����ωF���O�,2������ � (�=��P9w:�
��^Zi��%[8QO�}�<5�C�e�d�:�_�}���iR g� �׃vH�E����g��dL����u�`;b:� �{|vG�(�н�K a�L����?t��h���<�s���s��/����|����)��s5�B��W��.�[> �:�^�+�� E�=
�7rȨ%;Y��U|HDE��983'e�s����j����M%9���sN�#����i'ji!LӂT�1w�5�\�;g�yfQ�j��y�	;��~�P{fC�5ת=.GP_��5�~�Q���s�SN�`����U$��A��4
� N
'��F�q��ly�a�46���פ���~�������=��"��wz��4
����=e�I��*kC{s�����Yg��"[V[����)}0��m�`�Ԙ��n�b����� \<�����QW �>&�;&٣��r�	;_݈E��C��X�a怀Q��T�m�C�C�P�_�'s��v�ii�w��4����&���,���Y0V�b?���|���T� �H�BG� ϊ�8cpGa�r�GH�X�+"4��p���:�)�~P@x�����ҙeI���@��Ɔeնo8<��AX���(L�7�,K����1JĔ�C�`�rX����Z�ل�:�94���C������i�-d��oy�T�V��L3��)w�%X+��v �b�{^x�=�+���
zSP��3 �`,>��q�k=tt2i��7T��ھ. `>J��ޢ�K()�ό������<O����y���@X��,kS�$cO&{�a���V�I|̓Ї�9�<�$�9;[�-L����-���:\,n�Lt^x�����l->
���/JI��K ��C)�R���s�vl���t�<��O��]���eg����4М:�ZK��L����#���# �f��:�02�r��� ��G���W�)�Rv��,�.	 �zj�)�� �`�P�J@)�X��\��xY��öju׆�S�ʫP�����͢�O���J�I��;�*k(��������-��d('�&��i'C�ܩYϠ�JY:KgW�y����`0����"x0�m�k��[���~�Y�k��֣#gB�f��s�CPS"�%�N���;�$tg�q�:��clUa���w�+ic!'�AH��W_�q *�P�x�F����|� ý��k.�� ��Y`�V(�
CS vpK�=�Vj��<��������:�n�kL<7���w�(k6����^kΰ�4���*�m�i:��������H���@�@N=u�_ܯ)yL9&�]ך��\۵ȣ<`-�+O�(Aد�2��������F��)���:c`�e/!YDphq�-h\�-�/�z6քS�5��ɚ���kM�\k�I�x�n��~ޅ@b��Y~���х�ʅw��ShZ7!q?F�-T/�c���V��\Q��0T�g%��:�LXm�X�:�[ S�B1�Pn��h�\.�2,�S�V�d����"<�,�k��J��x��#��d"��)�
���kkY�������5;�nn�<9B�y1�=��|p_��lN@��Z!�٭�vj�e� u\��l:�R��_;OMݹ�N�n�u�ɱ�{�u��E�t���@��������r����5�">��н`jᙏHB	�ٚ�\��	�J9����hC��)� Kh����Gֵ�g;t�8��n�� ԭ�@�����T�� ̖��\s͛��	�����z�C���3�/Ą���k�-t�RL�C�Pj�'V�5�Ckx.��^;�����>Gy�X&\�T>{��W�� ����ڍ��U�L:��"���֥�n�^��r�C�j�C-��jEO��s���BdO�5�nv<_��:I��]{�o:�3v.����?����U��mj�\81���\�B��9���>t̡8�O�Av!@},�.�J��k���7� \*���U$���5��n��bq!yb1�8t̡8�O��Ɠ�������#� ����Aᕻ��2�:����l���2�����x\��C�j�C-���c)g.Ĥg#��ß;�r�� <��vk-!�.���5�!Mx)C�б�Z������n�Z�.�Z�Ơŀ}x�0C7I��_{�o\V9�舵;��35vA�'TMLZԂ�X3���D���d��nN�<�VP��UP�c�����	���-�U%I�|�z��}��Đ'�P\���L�ӱ9�%jf���ۻ�W�����Sx�f��y�����w�p�({��4�J;����u]�s���m�v;���<݁F/i�+����Z܇>���ؗ�Z$�����X��<%�h�������V8ǦiJ��篹�7.ktsk~pc�����6����ay�0����w	h�:;'(B�1��<��=kH���X�Ұd�i�p���� �G��8O�ε�����jd�a������S�49B���Q���I��2E��$J�����!lS��HR�}j�nֱ��:�¸P�(G�����*�	STM���+m��?�P�z�i���3�ɭ�.k��'�ND��Ͼ��|Ӳ��\�cۦ��q�AiF���3���yl5�ޥ�Q���\@W�Ȁ$����	�_����Tǆ)�4�R�<�&F����C��Ɂ0���r63.�䳁����ͬT} �0�N-c���Rjm7�	t�b��\��Z���|L����3��c�2�4�*L�Vv,��wҭ��®�WY�*��(�X5�9�td!/��|�6����иA(�!���~�0{�� <q�EY�VD���KYR����P��njS.��ԏ��7LcQ���q_�ܥ���k�K��򷵚u�
���TUb����m.���}���w��!����R��{������)�R�J8�BY��e�،,�pﱥ����X��݄�6`Nt��`57���X�Z���2a6V��v<P&���*�V���9,F��z/Q�)T$i�e�$�Q;�RQ0��ƠԢ ����UyOڳ�:[�eY�$��馛޼������9f���[�ugsa/e	�5��&\Mjv�	'y�3�+�h�Q���:p�S)e,yHm����:�i�IA �F����W\��Qb�F���O�a�}�3X~Q�	'�lZ�B�;�.!�����􋙨2�Y�a23�AX ���,Qas��i=�PLU����'��)|ń�
�<,��f-��+sB�E0lc��B�R��\����s�����t[=(�h\h�ƾ�����,p��z�v䡶�dRmH�ߜ/��a�����K.q�e)i�7�|�o-+����{��-mN"��f�3�4m{���/�~�g�����������F�K=8�9پ���x0X�W+KI��^��Wzaw�
�u��h��?��?�5!l^TB�^l��"�ʂ�	�Xf,p R45��-�P��<��� �S�Zf����*D�E�� I�~�U�:;Gk�w��$�¶�%2�(��%�} ��Rd�g�x�>v�ئ��`��!�9q�I��/��S�}˖-N� �b�c�	
�����n�+�qmI����R�禛n��e�ön�4؜��eq��5�v�e�k��ēO����η�Gn�X; ̍�TXj��P����#O�` �V&�����~�zc�e���0c���a0����9�r<�
����O�	=׽w�2Q�Ye�a��	���4������K���^ĀB=����c�'�"+�;�B@���b��H��ؖ���v�0�  aɀn���l�k(��K�K�'�`�<'8"�J�jW9� i��9��]��0hD[i�����Gb� �oj�K,�v	¿�� |�o^���M���Rl�C�ZGv�i��/�ܲvn<��x���29U�Rab�00d�*�.+<��/~�M/��<�����њ�~ɁƋ�n�wgl7�=��-e��e-N�(*�jgb��ahW/�ζ�8���Ga䅊sk[�wo�7��"�p_1���bcQ�����W���Q�Z�F�� ����9�m�v3"iv2��eIKܩX?_�I��g�1t�! L��"�0��7�W��fN!��ga�Ȭ ����Q�I[�I��֡���6\��5{�o���k1��"a�C;�l`�!��De�7��,���� �]t�c��,���.�j�	8H��l��?��[c��ҡ�<o�q|��7�������9/� y>��ڵ��K_�[�z����?��[������&+�#�ѓ���D������V/�3Iit��Fg�O9���/������c����ڹ�^���l7,Kؠ(�8�,ɫS'9N,�k�N�V��_�E��/F��,�V��hP��;)�^l���Y��>�������J�e��[�1ױѴ�Z���zll�iQ��r�FjOY���le688�+8���B�Q&S���;��X� �U̖��3������|��*}�]R�F��u�O9>�n��\�(��Śb5�0��{-{��?V��BKAE�`xX~�0m.F�lS�������}!?	�ɑ��o 5��O�=�k�����~�U<����E�����pa]*s.;���u�s��8������}C����|�+�|����d�&�gc4 T_�9�[q��
sN>�dg����q=��q��c��o�j�A��m��	;W��k��֝e�{��ܽ���~���*6�,�]���[f+���I�1!Y��h�dx(�>�����4 �\���x�w��M��{��^�A 4�Y8:"��͞�YO�~B�z6�h�������f��a��Z�����e6lY�kI\3��i�a�5��a�Yb�%Va�O���l�;.ge�b����Gj'��am�f�eyϰ�6sKz��m��3V�V��L-����me�ϵ�a�X��ڛ�u���y��Ō$7	D���x�ٖ��arL46�\�������w�f��ª�������Ҕ!&��K.�ĉ�fѣ?'�����I���/�r�s.s�c�$,��ER���/Ӿ[c^�G[0v���7� �@���`�� ��	�8�GO�,#k�~9W�5I"�"��M�[`�ӱC�g?�Y�GinEQԊ�x�7���SO=ud����6��8��<�ЦYk{��f`�����?m��v�~Ӧ'g|�L^�'l�':�	��ɁHs�I'������}��a�	X���Vt�� bP�����X��Ă�[y�jQ��<��x��8q�L:I(l�Z֞�a��ڶ�/����G�bGyӲxڢ�U���ȗ��;9�EHiɄ�J�;�K�]�YT+wp�,NSk�UK����F4dI��%�j��Q{�I��'��| �PA�.E�ȡ!�L:$MS�R%�cذa�O\,��ǒ�<�����k��a�/"�"�gԜa�/�C&.��s�)M�A��4a���:�|ļ��gø�a��Q����a�.spbΪ��	�L 9N}"�N?�tw�}���������5�\�D?c�FB��� �Cb�8�5H m#�!��̡{�<�c�����]�& |�5׼���~��e�y�sS�3����f�x��m�5f߸�߭VA̮�ꊼ�nv�VEn�P2�:O��@`�������?��yq ��
�x=�Cg3�B��x���0{�r׮7�*���XiIT)w��,�&�'��<֞s�����tݢ�bI��X\mZ�'���w�d�	}cP�� �Q,X9{����\��l��&����V����rа�9�k�������oج�Y� Xd,�tJ@�6�G�,Ą������A{k��<y�e"��_�җ<tJ`�6 �r�).p�o~��@g�}�?; Ä5��k@�� uM�����jC9 ��cN��\r�ƽ��Z �|G�N��W��Ua2��|��׿��w�
�q��	'�`�_~yg�^���9���'�"�n���e�6����9����	(�T;��L𓍇_��W��iG�{L��5��`�sЀ5Ƙ[�c�e��������V�Z�Ե�^�{�
�a�p�^q>�����Ͽ��z��y��=c��o��v\�E�C�����n'��X��:�,w�}�_p@�e aJ��c�a�p [@����$Q�\�.�b�f��Ȧ�Ik�T���m��
���X%���l������c�lz�NK'
�7A��,�iY�`Ū�Ŷ���<~�[�ю����۶�ڝc҈ݛ娋͢�5�A�6�o���-�eo͒��f�8lV3��C���x~&m*�!dG�i���g�s�1�MXk)�MLv �2�9�Iʀ���w0Pq��9��#�}^���o�������	�L�߹��s~@X���Ó�1��&���#X��� E�m�{X�|�V�d9���-&�pB���SR	�ym�� 2t LX�ĵ�8�3�]v�[ь�?��?��(9N>(�	��/~�k��E�v΃ �lն�Ap��6�m�G`Hj��ԧlb���J��'�s��o_V9^�{Ǧ���s�� c���^l�}�y����۶<�S�Z���+��C�0aq ����!�����eT�kݺu��7���$�$���4 �Xߩ pX��l²Jd�z�=�����ZOo��m�Ѵ�c�p�����Ǝ�Vi�]�h5'-%���e}+�ĖEm�-�=��� ��P�x� a�$��u�2��5sL�Ul:^a3=O����f��Y;^m֬����Ծ�w_qYFN-|b�1a&&�����ĵCY)���B��cp"-�ޘ��������W��c]ˮ�5���������7��#cx� ,тL���1��$'�m��r�s�m�	�9b�!�s>}���w+����˄�L��/���}z��9c��b���+�饗:s_�YI�	$M���h���cq��8H#��c�>>�<o�qr����o۰aÞ�X[���>y��G64��E&*��u���_d���o�O~��U��E�1�r��蚼2_���,ei|��4�-���%F������J�ַ��l���R#�CL�*+W|��
p-�Y�ֶ,�,�*����v�ŗ���g-��m0�a���,�u�ٞ]MU,��Fl�hOZ�3c����-�"l� ��ٝ� a�+�S�*�-ɩ��g�����E=6��ht����Y���hX-��*�c�6����_g���X�&�b�0Z;�-�`��F�H�?�2���!ib��hh�qMm)�?�'V�&�R���X��Zlh'_����Br����Tp b.(K�$�D�Lr_h)Ѿ�'��C�"�\���C��9�(��a��ǜ��"�@�`�,��]���Iý �<�^��Q�;�ڗş�Xg�{���CF�P��p�m߹C�ҵ�(���k������]Kc��ʇ�l^i�s	�":��O����W�w���>K[ W⃆���$E�<�< Ecȁ�g���̅�i0���I�~�s��f��s_:�L	9����5
 ��v �����s
�)���9b��N�O�g���X2�ǲ1<f�j�5�զ�oUb����q�2L��H���V8�J�!�'{��t�&z�x�{l��j���#,<����md���zWZ�ƶm�öi�-�Js��2���N�ðhO��2@��(�+�n��̄�[̈́T�<��O}JP��d���?}�R@�c�J�pѓ����R�,�қ5OȒ��EVćc`��0����&/?O� }�3oC�l    IDAT|�j�p��a���_��_qf/�<c0&�a�������>5�Y�9+�Ϲ9�p>bi�=��},�x�y�Ґ,­۷�5�$i%�ʧ����߾�䓗�	�����գ[nퟙ<��nX_������Wٖ����A��乯PԐ�a���D&l�N�� ^:�ق�K���t:�@��y0)^���q���| �55�+�eI�</��9�γ�/�Ģ���̢�n��X��n����{���VV��U��5,�N��a5��Z֎�;��!I�j�p�� �e���{F�<�i"��L���DGZ:t�eC�ۤYd5��j;vm��}�c>xh7M"9xfs̩M�,&#�KE1����4�n��IqL(h҇�-�&� +[I�|6'�OZ�9�&r��������=�dԢ���#�����R����ʜV"�/�*�G��:�#s&�~+*�>Ww{� �w�Gڡ|:��=��7֏�p�6�关��q� �w������cz3DNl��E/z�;���	<P;s/$v�`c��"cY�q�ߐF�S�Y>g����_�ӟ��M�L�m�I�r����v�o����G��:�Μ�8�U}+�5�y��+���g�j4Z�P�xb�$�j���x0Y���á�`��������x�
N�����c�G3ؔ%#`�SsLK3��YVi9�ҺmX��.��R�)�Jjq{��{,�����Z6�����*�%V�v:cV���ê�ͨQ������ a_�<��@���C����fU��W�Ht����[{�6c��y�؎];PX,�����^����!:�1x?X �-������\d!���A,	-��_AցE�,��O A��<���m�8�o �v��x���с������~�/H z@�����':��G���x���G?��Ge�2��_���:I@� 7�����d	@�R�3�����I!�$�3Y��8N6�|�o]�d@xŎ��4��#�VWM{���8�t��o����5� ,�S���LQ�w��*i�����/ o�V8��I"a �)���/t3X�k� 7��!��{��k�P���t'-���ε�/��(Z�T2��^�w[4z��'�u&� �V���X;�*@xM͢����aq5�v	��Q�`����펼*���DByP�ØV���Z��K�i����Q�,J|�	�s�T�ik@�I:��B5���̈́+z�@�����2�q�2a`8|��$�[lsR����
��b�k�qA*��s ��b�1�áDԊ<�rl��cɄCfͽu3aƗ�Z�Ҧ��7��1�7n��G;]u�U��}���Xrh ���'���'|&'��QV���NEf���yqέ��Z�ǝ]N�8�6���w^��������j��;o�=�R�#�Fn�x����r��{k��ۿc{��u�T��<�FiHҠ��cN|�;���d^�9A#6��/��l����'��AJ�22�^ �=�q��(`^;����n�;�.-A8F1Ha»-�{��L�rĄYҮX-��c�%�yâZD?��@�9Ⱥ�� �Y+�!�c.+�
��ؒw�5�NV�H�p6�D�]{v;v��qhƲ�	�	��e�jA{����-
c��o��+�`EL�4j�έ��q  YʄY걡�p+�S�E���X�򗐀�sa��_���X�ɯ盭m�N?/9B�7�q� �u�n��O���6,�$0��?�tX+�p�X����q��״��44?���tb�C_@���/��R�7iǟ���w��noodsc�<@���e�{7<�l���n����L1xJ�`Ő�%�=7Xw�q^ד�)�ê"ݏ��Ӈ?�Y�t�M�'�h�l�'g _��>�B�T�%B��l(����S�f�����B��jn��a�#��,۽���أ#`�E%Nz� Ѱ
L8M]�)4�"Y�x�Cj0����d�I9��������׃ӡg�4 l5��9��>�яt������t>��оfa�c�	˯�s�Q��I$����d�md<���BR	��c	�|� J���XwH�[�O?��uc*S����Eb���ǚ	�ϸ�L������w�	kH�j�P��i+B\�z/�g�+	��"��t/�"p�9VQ"�M�0�JQRT9�r��]{���}��q��y���Q���P�jN3���U���/�c��ۻw�'+��t`~j��0����d��<���48C� F������Tx	�F�����A<���`Z��c��#�~~5�ن��y(�9@8j�#��{��=�-3���,A����6c+V�XқZ�Z�	�{Z2�C�ps����,f�T�פ��4�Y#^i{��>��Ԧ��1%�k�}���T�͹Js1a@9��	?� ̽�AĠ'.���������cG�C��c`���`�9�T��}|��G�3�I8�]8� a�5!�<�����_�LD%�������!��� bƳkLз|/Y� #sN�j�n k�L�B!���q"|�aI�\�q���u�D��Dj���y�F�����~k�Ax՞�n�Z�o�Y�*_�o�y��G�e�\nO}��;&<������(�a�_q�����XB�-��D�������;5�u�D�|�΄��S��>�U�2�(����b� �ǹE0�ֈ�,Ax`�f��[2n�kWc���ZeƆ��&��N����v�.�o=羞�QTS#"���URSw	WJM�hOk�LM��Շ>��t�9��҄CGR8�5��ßgt����,�)�i�L�C,1$
�0�1@VĠ���9� 	�Ysį��x.2�p��_p����/�Y]�7>X�9�[��$k��m�I{i�S,�p�=�UD6�X�)�X�)�_�D�(� ���H��e�b���gL%I�믿�ͧ�vZ�f��W.B���?3���6��!k����#���ϿЫ�T�&	Ńk�X�y`�[<�8�4�@�QQvV:�A�7�/`��8��C�r����}��sˑ����9b�q�!e0W�#.��b7�Jdyk�V$;�2r��>`�.�plQV�V%����:m+�L�A&L�Kg�D�)mY@[�����F%6�䊈	��	Q��m$:ڲAs'�t6XD]X�Μ}�`�s9$�c�b����v�-Ą�cN��B��h�D_�rR�����B�L=͇n=u!Ki��h���}bZ�З��u2��C�gZ$�Gat�Ƶȅ���d�z���&|�SV��WI�q��9a���r��>�`҄2L� Ua�*����5�/�o��^K�\ߛ$��������SNپ�q� ÄZS�Z�EloT�F���N��Xjδl��՝���Nx34�J#�aa-���.�ք'U�X��Z�X͘��A�j*�.!}�L8�T-w/<�#S�p�:���+<�"�T��{lE���?���,ߵ�*�5/{�&�5r�iZ�cվ��6eq�>w��Җ�+�sA��je��q\��OY��cʆlĞb6|���������d������G?�1DZ�d��jr�=4i�R���sK�q:<<f���Xf�&�)m��	� e*�1�m�p�R3��g�1ǘ����l8)�pqYʄY�cgc�ZS��-+�]�q��r̅���sR>�;��?m���e�"�[9k�gQ�V���\EbѶS�1�P{�f��o�qE��0[,&$Q�^�B �(�`�~`A��$�Y��9�ƊA��P�?n�⁤�J4g���r6h@i i ���x脜�/%L$��#�4�(���iIԴ���%�\ayT�(�ytĊ������F�|�KƫV�H�Ȭ�p�C�*}��(�S�"G[^��K[�E�(k\�#��&Q$8Sʒz*�3���3,>�Z}'8[Y�~ddrY@�I���c�Q�θO0 ���zʹ�@�u�j�Q	a�j�j�9M�p⨏%K�\_s,�� ����{����\�x�ɿ\�/'��_��x
�R���n܇�Q���e���A���b�b�ݖ ��/�
#���f9ڰ���-�p��И�Y��H��2�3����2���~�-��/��/����u�-���	�\c�2�wZI�h�������Ԑ���JիÀT!l��,J�Q�7��}V�����l�����c@���V&�,��c�}�l�N�Ɖ����0��,A�m�h�ab�Ҕyw��>\�1��uΫ�!�"��|���3,[>ѦmЬҶ<�ld�1a&��61dEcU�"\h{+����<�ؔ���K�FAh:s]9ESE�/���1�!�-3�X�/��J�S,5��D���̧��a�@�9����zDu&�8�� _��cT֡p!|v���/��4~��y�RP}�ꫯ~���)���d����<�4�pjUY�����%J�����>���2�H9v� lYW-&D-�a�L���"D-�A��ȧ-�4l�0�p� Wr��,�Ȏ+�E˨A�����Sт���F�ϩ���^{�e+N�f߉6� �~��ޑ�b¬����M�y'����j cn�?Ŵ���9� �|���2���=F�_�R�Z��.�*G�sD ��e��|�X��
L����+��\[	�}��jĜ�[���	/�8�!�MC��M��h,�3�|�mY�a�yI��tssi�����v����F�đ�NTCΦ	k%�3��.�@���>$I�˄�j�~h"9� �K/�ܓ!�J��ֈ��wX4r������[gUK) ��XTi� L�ܴ���R@�eׅzV�q&iCr��QA�cW\`�$ =Ͳ�S����0���yj���oM&�IF�$t2���>X�ژ��!kcV�_&��JJç_ m�C%� F�T(1i��g��Q�D���	/��1�YHHr^��#Nrڗ>�?#�x����A����1"���>d���"�K�-/dg;&���tȴ�H�� �CK�G�<z-(:����&_z�;����g���W"��	��6�&�Tc���� �!�sp���39��%GT]�hg0��ˊ�JdI9b�%#�Z������'2KҚeq�Y�� �#T�_���˗6��w6�$�W�k�gЩ��d���FO�lų��m� �,�ѽ{��f���^�2�F�T{j�G���)9�|E�p����`�&6!�h� �����7�^�0a?���>Iԑ�|���x�\�+���0a�@E�f tZ�	i�(���8"p��
�|���x��F��6n�ܦϥ�ӧH�:Sd��R���$-��]J_���l�fr�"fb�]-�"�)ZV[qLX$ܢMU0���f�{m�j?�Q��kU	�y��р�*�P�;�,11�Q���B :"�+%gv��뼞0�I%�>+���z��l�6�ɖUҊ��m�M�jᘫ�1iqMv[TM+��[��Ow�#.�Kf�;YSLq�&�a�c,_y������h��fY��Q@���̈́e�2Y����U���r�i��M�|���5�b�3i�Ì�WIH Oz��)r  `X8p�!�(*JYv;�y��(�N��@����!X`�B`����I�� QO�0���F3>�Ѩ���o�)���`GG,��"',V�~�n��cDFĞ�\Z��`�>�/_}�տ�sg��u5��թ[��i���!u�:�������D���`��SO��CmR�G�����.����]���c[,ݽ�l��!jq^5j-��=V#m9���kl Zh�*a��j�o���L�D̡^���m��\0e���h�'Z��X���Q�3��>����4X%�҃Bט�r|Jv�x&.Z;(8^+�ˎXv�Ez�yU��3R���1�n���:Ąa�%bQdn E��`� ���N�d�J^�| Y���IW�{J�R�������S���g���.�Wu;5�ĈC|���*`�v�q^����C��F�`�c���}q�u�V��&�LZ�S����aM g�e�p]S��YAè�j���|v ���m|z�*=��f�%qfg�;�֟��B���6PkXOk���wZ��Vk�|��vj=l5?M��*=��V�ޟ[�PԽ�l7.����
�}#ϝ+I�>���~��UkE+m�~���Zk՟b�jeв��G?���zM��[�_��~�U\���M:Ҡ�6���H�..���Ċò��$�����������c.�ﰟ�]
�׸�<~��)r!F�x�<dRr|jQ�I;�a����J7�}��-����B������=Q1�$%-���{~�%�cMDI�����g�kt��>�YdOq3ܛ�l�w�Eڂ�BB�=��Ӓ��x�oX�d���4Ԟq���nMb���g�S@��0Uוϙ�ܸ�e���A\#��al����X�a����^22'.��g�L����f$��@�������ZW�hU��b��"�!�	�[���ZwHXk�U�j���T��ֺ#n,!�(��v��������͏;s���0A�>�<�ν����y��|��}�{�ѓ�jé6<���+͟�gޞW���J�f�ғ?2�������4t�})�R����fͭ��Y�)U�2���Ŏ��O��;͍.a.�p��G�s�A�[ޏTSo�i`d��뻺ӷ~�5���z�>4+oo�?0��fW�wݞ��pΧn�b�A����ٌ�Dd��@ϧ�R����ar �5�/R>s@ǙT�d��B:K�C����&N��O�y�:���s1�`��1�J�@X������0�H��m� `��;֔���˾k�5LG]���0<�L<rue�jo
ޭ�8+�3 �A9�� |�����-����h���8k�O�B5�.� ��wDo
���W�s�_5�5���R�|�Bc5>!����T��I��q@`7�����Cs����ݝ���Ҳ�H�<|ߔ�ߛ��G<YB�!
����9]����b1Fa T�h��l�+q��k:X�\�J��4R�3m������Mw����4�wn���<��I�Q�� ����YC9n2�e����HhG���mTpqq�!m�̲��g2cLؕN���;qO����xV�F�q5�u,�8(f[��j��X����`A�v�(Q�6����x�5�hg�qħRg���{%�8��?JأP�K��w�H'���1w����Q&��'�y3�ޡ	+�\\P�a�N/bt�9�����gܪ�q����1A8�Sȫt��z-k��*}i�V�	�{�7�=u�t�K�z��<�r��Й�׺rv}v���~�#�d�����0[�0.rDd�ݨî��H��oY�(r���M��J��3+�5��`eϼ�ܬ��42ܕzq*��	��;��ul;D`G������y���'׍S:�����ц�e9��x�x?l�)5�F�|����e;D�}�m�q��� %��I�siyd��c�D;����+��}G ��y����Ĉ�v�s��&��vm��x���0ʛ�m0JL>�q���:����3����4ox�ɀ0�0;k�	Ä��p�O;�y���J��p1���r�Ƒ�ϲ G%��wݑۥ�+˶L� ~��s�B��,Fm���C�eO�>�����Z���	*Sw_ޝch�Z=/ި�i��)'ú&\�z�����	�yϏTEbIi`h0�V� y,�����ޑ�T�w��=�RmhG�&�N=�p��:C��� ,��ь�6|Ɏ�%�C���dJ���#(	XN!a�q#˩v��:_)I���"HH$�t:j�x#��b�`Tn�g@��8˱�c[ęQ��9�_���t�o�{�A][�;,'��4ͥr���qF�����ׯ?���,:�m݂&��2תEn�rr ��I��ȍ��J�NI�C�C��	�����F�GϽz�w�0�#�E��0�X�Z-��HwW��3�D���ONVv�����W��9�C��v�V�'��x+���H�N��ùJ��m    IDAT�r�E<p��Q�w�``뮧
@?RO}LS=�{G�}��4������ԗ�#�4<8��K}�l4�8��٥��LB���k�Q�ߨ;�3؟�E��i���kp�ZN�}6ʍ�ow��S5`m[���R81,�6�2M���(�U������	�n�1��o,�1�Y�`�-r�a�ܡ�R�Xvن<�P4%1��` g{5�0�I��� �c �V�����	FA���W�[����a��{��-7]6���ı@�o�G�$��RHC������O������
�����n�ǘ{�D�q�T5=�c�
��@h �f�uో\�Y�������Z����,��\�I�������`���2-'>���`��]����袌"�ew���ݬLN�Yը���]i�p�W�){�9���T�	�y9��3E�����4_s��؉4���O4����S:�:8���I|ﾲAX��Fg4�Eu�������v1����m�]��x Xx%)�7�x�V�C���f�Q��Ⱥc�&[�c1me�Y6:g�D��O����a N�û��㽭�Z�FR�O�]����not�)o|̂[}ټၣ��#�,MG�<O{`�,�t)0@L�#��,����H����F� ك�կ~uf�9²��_�%}����F�lC��:t\l0�����@�DO7aa���RO_5m��K�>��ޮB��W
�2�YlW^��f��sNI9�0����bۣ"�;�,3Lf�gw�kp�t���*��ix`8�)���]��h��3Ə�k QFh�c�'W�;DD�O��9U�N�DԣǺo�X˯3���d��8/- ���h)A"z�%b���l���9^�ԁz,`�H}4c�9?ړ��l��J�2�";��C`x�@\߈+���X2L���$�'F]���稍�GA�̎���3�}�­7_6����f���������@魥�G��z���ܹ{��}�ĎJ�!���cB� 8a���I@dtTSw�[������8 ����,6d�Ҙ��[��e 娅��JA���ʷ��b��w(ݦ ���FW�!d�P���G&��.'|gq�+��n�1�sfj`���8#V��oH��t�Ȍ�-��/�F8P�q�gnԈ� �0Y��y����q222R�V�W�^����������qo��eF�����>�ꛛ����%��}.�g�����<3Z ��;zEu鄃�`h2 7	?H�c�Q�6��F$������Pl�Ɉ��h��2��t|���f6S������j@)�߉�!18@�~&���0�S��3���v�Q��0��7�*gI�3GI$��N�Wv�t�pT��U��O�Y��� |���{���n�t�T[>8ԟ*�=iN����כ�?���'<6���?L7�pS~xG&
�X�W��2��T�ёyg��I�u��(lEr�gf����hv��yի^�+��@�0vT<��L�����=k �����/��>�����ӟ�tƒ�N;-�ڏ}�c�8i��'P�p�	YZ��%��o����p���*P�o�t_&<��U*��֬Y���2a@x��o�t��m˙2�T����ZZ�|Yz����n�rC����#�2Y�:#�9�@N [�8!��lO�6��xE��9�5�C�1B>�y��K:/���V��{�}��5S�����V5 ��߮]�6˖��H(Dn����gdݖ���o�L\b��g>��!���Ȑ�W�z��椁�q-�y3 PwvF�X�j���޹��9��d�	���+_yR���M_��������<t�=��fu9�0�0
�;R@�'��e:�ta� ����f$#/8�{���8H��V=��L����Y�k�o�ƍ9���?������s�T�d��ߌp@�$�j�9���~��8j���c�0��Db!��?��$����3�Wz���z}���s�ʋ.:�裏�c"�9��Fh���vå��+�g����:��?O��vk���'��0� -q�)����lt_""m[��]ՠ��b�w[#7�|]2��f�੠�,6.��d��D*v�ؙ����� }��~�Yge�ǌ�+_�J��t�Iy{�ؗ�����~p�햸; �n�`~#���J S@��	�u$�Fd�w�'�
}�=ц��ow1�p��犕o��G�a^t+ <�"�k�w�#Z�^�����~�����s�c3� � �a6�y�o��%nh��~�s�˕�s���>7ꄓ2�u�ע!�hB��͵�1�i�0s������	�N=���p�%�4��������H� "���,�e��A3k�M+k"}�S�p�br� �W\qE�>�ឞ��^|�9aC�fo�gEo_5uwU�҃O/|����?��t�/�z�}�
�ٳ�l�~�2@�QG����k�"F/�7�q%
�d���'���m�љy��)���vr/�s��㙹�L����k��f��0�8q�� ��_�H ]�3��
p� +�~�QGe�fd�=@��dʞK@ 8�}�o����+�+֯[wnGW̱Xc��o�l������R�қ���)�9�yv���+;���B~ (M�e��Z����<������+���Y��-�tR��Db�Y0�py'ͭ����L�&w��؀+4[�4�+O�r �剋����&w���fj`�5�bR'���$�����~&h��)�a�G� 4Y��~����Z��֍�pI7�s�x��g~��[2^�j���+6���Yf��n�l~}��=��'�bɲt�q�������0�,a m�/�1!F�&L��f5���e�\�E�`ʡW�� Yco���Lu�Nfq��IE�+��d���yqE���������@���g����]Q�#��������P15Z�hq��C� +�lGb{��h����a���+s_��/��8�8�.�i�;�w�i��V*�׬^s^g�#N;瀇ܺu��{�Ȋ���i�cN'��������?�M{Ι�����a��v|+���n�v������O~2��6c�,��F$e�mres'�s��
�h���I���,Nڽ�T����u�KY16�nq��<�{Ϝ;SS���J,0��MDF�Y��=&�r��/� 4�4\���0�p�o�;���D]�w�e��&������^A�V�t_�f՚s:
¤�|ح[7Ww�Є�ki���N:���Gw��7�=�Tzs�'t���&Y�s#���k|!�Þ��?�3�ۿ�[�B ��s��:(k8� F�1`׀.e� e�;�	�G��Bx>���j��:�����['N��aДGО�#vU��\�� ��^t�EY����?�#�d����?���o0�Q b��׾6�� ��nr�{��9���H$Տ�vf��)��ȘE��QЮuww]�~��7tT&����o��{��O�ф�Y��c��yp����t�w���"��K��� OY+� A��d��J�2�&¡�4�!`�nXhs�4䪫�ʂ��J���54f hW��PN��N��v���� >S�������������vjv�]Y0^�[VŲ�����l�1c�g�}v�	�����Fg�`;��&�� ��A	��s b���I�93(�b�.�Q��bnÆgw4�;�Ϳ��s��S�v�sC���_�����$n^�|���
Q(u�Ȯ���p<������ׄ�?�ъQ��/̕�bt^� �ד��f�\	CÙpyW3�VH���it��1���u&�{̲�5�z�_��;`\^54�	O��g��d�G 
o�۳�K�6������R�>��<�Ɩe�XDz��$n �a����q�]�'�;,��C̈́�%��G��q���wt{�%����o�_�JN-�F�J�?���)G�'�����~�n�qK�XP��S��0.� ��̱_#�3� \��9DE�(X�3�1�?'��	9do�����a��"G��-o,�I�mv���D��`���@t�KYC��e���L�`�Vlذ!K���Ӻ�;F��ۿ���س)���! ( 6�G��G紤���lj�#G
������>s����y��כ�=�,jh��g�K۶ݗ�~��t�I/O{�~��~��F!e�N	F�_�# ��K:K����_�r��-�y�a�/x�r���5k�Ne��LN<��� �o�FFD0�.ӦL�>��g���ەe�i�d�Tˍ ����͙����Uf��n(��L]���`R&'��7~��,`��'V�� 1��b�[臨�p.�{ Q��#����(�����ի�\�b��v����]�����7e9��-��3��N��f��K�����G�I}�~���0��.tH�V�e)!���qn�"�������z0Ss
��%q�X 6���#x�r:$y~�ɑ�ӌ�q0������kT��1F�-����5���
����=^Wϲﭞo"���xl9,��R��~��(�Y�гo䑳��F���{�R �v1f<ΞʳJ�#H��m�M"��%쬁4qd�da��^�)���8��� *)FGv�Z�z�ʕ� ��nټ��}�u�����#��?-YrDη�*5m5��Ί
�~K�(}�m7�V��^���F�wݷ��T������Z���t�TA�rǎZ�.Q'�Af���!vJG�<��&�',؄�+!ŭ���k��xJ����ࢮ6è[[����8��Ȩ_��ٞv����a�!�dL��nx�mI��6NV�QB�OJ�F�����$���	[X� ��.���?���!��f�h�h��F��.ᅷlټ���c���]��7¦��4��������ex yHqTعy�^m�(�Ȥb��=���P1�Л�q�2Io�6IT6��ow0���pd�J�*x���A�E0��z.l��L�S��1F��-��'	S:;*���L$�re3Ze�����|Yg?��>��ːe_q`��9 ��Vl�����,��
�'���q�v�ߝ��g��]�������h6�C��|����E��o��	Q[x�-���C*���Hv�U*�y{��jW�>��R��E?!�������Kv+iTP��9��ў�q�^+�����Kc廨�L��L�}��F�)�O��m_|n;��c,c�0{����k�S+CZ�aꋲ.�tNɇ6a��3Jmۖ���3r��V'����2U�Ҏ_f��]<�w#����A�ߔ�l/�]�����S��о֭����)H&�G��ܡ3�BWRg{Q�Q��l>�jժ3:�	��޼i�4�CԈ���P��+�y�{k�l���
��x��70�w
^��G�|���]��q^�{E��4��=;�Qv�^\�5c�.q�ȭC�7"�����ĥ�tv��#�N�G:A�rQkC�f���#{��Ap:۾�{��r�38I����?���U�5/�}N-Y�ٶ�ɸ��rRԊ��(��ygJ�_�g��c�?S�֫�R��D2��,�D$���J��yΎ��[6�ڞ�p��I�ၴ=��k��OIc�Ԝ�8*;hQ�N�Ai�\S/��0��זEG`�#�*ǎ�N�@�B.�� �p3:��Og�dY�I&�(�jL��п�y������~G��҉��`��N�M�{J:t�Z��$5��Q7XW��������՚�f5�2�*)	��a����˱�M��Hg�;�	��y�������@x��n!w�15�UO��	���L8�q����O�n��4����5Em3o��:�h���ָ��8�
�ց�6�8pJ���{ �a��>��G��� ��.f�����	�'L ��� z���Q����v�{�ʜ�҇�oY�ˀ mI�	��� Sf�T�s��>��������Y�ǎ\�GR�wfBq�Jh)�%�ҁywg0�팜:�e�\g�b�����,������R���U�N�a�ڞ�ێ��Ɏ9�-��	�h��6,&��,I#��� !�Ƒ:N)��N:�1�?Fi����S��`t*HG"� ̋�ynS|�8�!lQ9��Y6��g=+k��I%�&uFAX=��pʱ��N$�)��κ0�[��e�W2 J���?=�����G�đJh&Z%[��,D`�5�g�����Z��c���S��T��0��ݩ#R�������X��uhc���|NyIሳJIbw�g�$1���sٯ��R������Z�~n�ʕ���7�ߐ#p�EM�|�lo4�+�k��>t�si�udgN�v�!��=Ǻ� [�3Q$n���;K��q�-��]�/����A\ո(&L�PLØ�u �h�>#I���eS�9"o�z�U�]7��8c�{�'rvz���������%3b��SN������75�K�_���e��o~s[^d#�"	�7� 6��~X��C�^p���X*�c�2��h��I'�@rg��g<�`Vf���vlD"!��>�6���[��OG��U0�@�ddƞ�3�,����V�^=} �(:�*v�8-K�h�3���\�� 0�����j����@
`	[24�����v��rm3�3	�x)FX��&d��> �&�S�k�0a�2jSiߩ���p~��|֡e��$a�h��?;ǰ��$A9L�A�#�Hc� [����`�.�k�\���xΣ=a��S�^�}h{ڗ�|�0�^�r�=ǐ��킢��l�ϱQ,��V}��~����ҁA����l6bV�Si�f��e����իW�:mL��
��-m���:[�L8���P��u���a�9�IX���z0 ������d(LU�6�9:*�ҹC;q䍨r�B�AnP^���7\[�w=�s�<e��� S��v����ߣגf�J��A� I�=�i���h����m~Е9����r-]~�3�%�����n�àMx"�Jy�=8�<����L���9���� 2�2�;x5g�o����,"�h�e�Fn�Kwww�A8�	�~��yC�O6:b,9����� qA�U#8����\!��P�*6B+&���Q^�̹���	�+�|yǠ	�1 c��YB�Ш�{����q a�q�kP�g̯@�W]	�DD����Sov���:�6�kE���I=�qw���EG��Xe���}۔��3 /�~�����3�5ϋ���V��
�9β웂0ύ�20�~?Q�PD[�n� �#����s<�Y�/�p3v@��rI�m�i���O���'�v�~q����oy ���*�,NכU\������@/w�����l��tZ-/?�n���~�ba6����Ɂ�@�5�N���AE9�c����܁t��=\�)@������O[I��TR��xw� �m���$�h�q���b���؆�q���oAK-U�Zߋ�t�ǁA��;�C��bߚ.K��-Gr6D��3;�)Y��r��>��������_|�i΢v����qæy��O���}F�q��fc5c�>���]��@��)_�ȷ*�n��ǁ��bGta�L��b4�XSFt?e@�Fa���D��q�n>˰"s��щ��g;gy���;�d������:���d�N�e�����`���]�F=��D�1��vv�qê<��8+⻸�7��LT0���#���a����P�Ѫ��V<>2kYh�-b��e��s�7�'~�Z�Hi�	��&|�ƍO�hRw6�\��f����@��M.�"D��м�HV���)T��+O#�M��݊I�j��{3@m��~�!�r5�������}���L�-�h�YM����0��b�ttbK��[Z�N�k��5T�G�=ֽ�S
�D@�H;�>�0m�2X�����]��\�/PF����w�j�\י�������ϙ��Ug0�%�����=Nn�k    IDAT�˃4��Y��"�Ł���@O=(��V��2�6�y�#&�Z�8j�J{�E$�M@x�T�6l8�� ���s�ϖ-�������Ã�T��Ô AB��s��E��e�cQ}��Z� ���S�����"��G��x�؋����	s0ؘ��%�t^�&E=��3�Y����&�-���=��*I����M�������E0�Q3L����zR���U�V�߸�	��d�q���UG�{��j��G�$c4���pu`y/��t�U@�r�dAXP4N�ε]`�w���l�W�tf�5�_�ڙE���c�g� Bd��PgQV��������������s���?��-�����"�����ܞ=ROO5�n���7�7!G,\�o"'3��놝�)5H2e2��a���9u4�3��!5 8�xVxq/��˼;��G��`�>\d���
�W����FA"{�f�jO��k45�hxh��>u�P��������G�Y�L�����APo0Z��9c���(/�e�갲R�h���9�&S�>���;�G�)�DBP�=p�	^���:�̤�}�M#A��z��.3β�j{�g���@}�x�xԩ9���I��a��=���l�H*��%: Z�>��o;]s�5��2(��� B�����3��DT8�44���^,V©N��"���y�Z�>
�gv�;���������I�#��R��''�a�2��k#�i����'=�������
��蘌^T&�H��*/=�N��n�R��SO͙�	��J��\���.��q=;�#����jw�N���-�>RhIN�uVݷ� AxpT
�1ֆ��p����k��f�ޣu@i���Z�:.ue�.��Da��brωr��Q��q��q��u1­�b�AX-���]���h�/�}��
^��"(:+��	�Ԗ������@��B����#N��lZ���S�X'�����@�5V�Z��г��5�yM^<"	S�i��#yP���0K��4��[���wY��XZ��KRJ$�v���C�$�[B������n�|����f�\��g�s�q�\Cs�[jw�"4����?�fAt���gW<iߘvqϬE&��<��('��Â4���"B�Y��#o�02Ȕ|.='�(��]5�I��J��n�E+Р�˿� �IK	E����!E���s]ų\�&�}Gu��q��|W�6��a���;��&�Wgk���=��C��S�B2����燫�U��+���t���SdZV`�l�O�}���$E;߯�SA�A!�gGi���f^��G�AEY]B�8���w�Z����6���;V���@����pҧ��ȭE=Iۍ��;d�1���	\�E
o������.��]_��ɾT���᯻x^��ԽO��@�1��<�n�����xĥ�D��k�ߴ6+���,���@�a�8��7�4Qf[��|~x�J�2���e �4�g��ѩ�]g[Z����K܅��C�A��W���'[�� \e��@��G��r?Ti��~�D�;[�ǆ�|�̻��	�!�L��m<���P,�ǈt⺪u�_t�D|�d�>���[M���@g`;�/U�:���6�zs������z�r#K���cq(���`p5jG[�
HJTS����b�z�$%��-4��6t��J�������#�m���
������B��5�C!��A���2-D�V	��/��߯q�0Wo7*"����?r�oi|��x0l�����v+g����gd�0�E5.�(�U�Y��6A�z���卣��pBq�[�eF4Q�Kv[Un�D8�;T �����,�X Ti!�#HZ�&,�K�<�u0J"���K�� c�v�!����y��!E��W�m��|5mA�𝌸Z]}ʺ*1~b Q��	�Sv�]�F%�Ҩ4���/�q ��R�8
��Al�M�#�7a���0�Ã�ɑ�>�+~���~�0�����������9���i�<dF|�)c��R���f����s��q���G$־�ݙD%!I�l�or�&b��i-9��D��?�{����I8]�����h�&�H?������ 4c��~��j`壬����+Yݴ��z�lL	8|�SLT��}�'���H��������9|V����鳯L�! ��{��������Mϡ`
*�e��V$8�O7�=�g=3W;���Q�M���3��o�R�,�>p�;�xS*��g�^�j�g?���ѹϰ�0�ik���O��p����]��f�V�ǃU��'sD���{�=����Ue�±���-�2{�^H��� ۆo[���m�����+�_��EAA^�U
�����!(ĿBӯF@^��?*��紉�P��:)��/�� ~����n���N����öQ�*�H�_F��}��!,���bw��Wۖy��}deQ��\C�`h��(���+���_l�N8w�Sد��E�6��%�6�e�§#���_K��R�v�O|��Or�?���7�-�a�*�z<GĹ |�BL3��D���c[��0�u��#�������!2��J�G{\\\GYY�ί�.�
T>}�lE�F�Iʷ?�M�N�o������$���ةA��E�f;��L)Y�O�a9�6}w�,��on#�\�P���;P���x�����/�u;O��ZC}�&�~�������;ym=YHZU@
��y���NOG���2: ���̴}�v�6��7���"d�(#���h�&Z0)�X�_��v|؄�N���|q0�T�P���A'`��0z_Sɻ�X���C�f�m�����
Y븀<��̠n���t%�	���d�A���)/ e
�US��������nMYz��v���Zf�D���s �*p܆�n��]�N��p<��� �����]�Y16�OpQ���.OIl�sM����п=7R����g�iv.�o����}b�gr��M����>��C�i�mq��6�: "�ɢM�jVH��,�}&�f�H��	U���q�]-���͉��70s8�%�dq�+ű�j�XY�x/��5m��;�����8���������?��B�ѝأ�yI����"�m�y�r{G{�?A��N��}��^3eR��"q�(t���?hP�U��a�&Q#3Ħ���E�nN�x��'v�&U�۬#W�Ϧ�\o�sa(�k�Gh�O�T�QWS2�Eb�zB��c#��$C/����(�v=v=9���u�Z1���G�Znj�G\�Yp΁��wT��U�H���:�#�BP̟����C�D�����u�׿v9���F��G�U x���HV���j\WM��a�-��G�I��Ԙ��-m��/m���UP0v�,z��>a^��Ⱦ�z?ز��S��e��Ci�ĜK�4p%]�N!�d�Ϩ�BW ��k�����(_�V3G܄)��5�Yj���!�b|"ѳ#���UTTދ1��r��2��kP��N�i޾�$�I��^�A좰�.rf��`��8i�*!0�y�?X|q��6�IɲV3��{��O�������y���x�Y%���=����FoZd?K�~��
�����C�����{A~+���5ӂRw�ٸ*�F�o4�7'�{ �{�N���Y����O�4D�^��c�y���"�Ju9%W��ra)��]2���z�!��D��Я0���<�x-�ݷ
�3zܐ|����Wh�x��\����D���J��AyEx�1@�(�q�c�1�C�[!V OK �C���*����P��И���z�� >.�ht��R���%^�@ no >LE%��d��wx��<�)N�y�04>®�|q..E�I*6`�����(�Z��^k����w:�Yج�o���KF��-���GP�X�uM�c����39@b�����=��� ~M��G3�l�?�
JX����"��5��ʡ�w�vC�&!�2��Yu�����wһ���j�ޥMoy�/�� O*J��ts�x^���(l�������k���.��������Z�ގ���M�%4�3�p�+����c����}��8�����µ������l�q����Y#�z�X�������T6��1S�������g^�u��j״�a�_i2�5&Ry b8�?���i���QLݡqn	D�/mZ&�3eS�zJ������;7�<x�N4�Bj�b�w����|
`�Y򐆈~�!T{�i��{��]D��.ɼɹ�zZ+���!�"aJfQ�}��/Gc�lAP����Fc��%���y�ڀ�����ii��l�7���SE��;T��Z��N��p_ޟC����x�hg���J��m٥�;�qr�R��e-%���xO�Y17"h\�F&����:�.yT�?���Я-�K�S��'�7��
 PQ����#�Ty�9���5PJ(� �TF�����F{p���x���M�[D37~�i&��'��Mrnʫ�v��B��7I��c�ޒ���_����j��j��F����}1�`�x�'�v8W>��j���2F�?
����
FR���h;bo3ڀ ���wjh�m@�yS��qV�k�;��2�m��1���W1�p�����7�����8�K�۴���&�O6�/��h�f�����<����}Np��N�yh���9~7
y�nM��.��K4�Cc��_F��Å;���(*m�^|�}���2��;A>Ç�,�t�a�s�WD�EB<�� $�(��^c2lyD��5�U�5��fW y���"�quޯ�+s<���A/W��֝��3ٔ�5���p��Ev�ߌ�^�TD�-&=��+%"�k..�Q{/��B�� .	���"��˰�D�һ5�W�1��Bbn��u���{X���rD��o$�t64I
�pV
5��ж���Ñb�
�_��'}�vd_��2��|<S�Bg��>�HV#���4�v"s2�g}�xu���Q�,;+�<5X����ż-2�* �jܒ�Xy�zff�v�v.B�>��3Z�}o{���*��8�z���eі��ڙ՗[��8�h��	@�@� ЙI]]�!�����A�g޽�c��#����#����z���VBՒ��]h�n��//��	>7�+(w6���ƣACcu$'=j��V0����&��'Q��)��"��6��0XP����D{��ǤrQ���QX��n��g����e�{%`?<+E�	������ID.+D�,d���պ�TF�^L~�^~�A��^�#�^=ZV�	O��pS�=j�DF���-�1X�H�I����#�W��PS1�����z��.��a�a]u�h�@���;i�.P�<Rx�>c�<rr���19EGu�l��X:Q�d���� ��'�Z��t�g��'1��?.T<��X�V��T&&�2�t����?W��kȬ܈�K�n�S�;y��>N�%��R�N�[�eL&�|�H�O���{�t�D�h��H��wyZ�6���T�)l8e�ǭ�v�ʂA|�&���Do@0�juʠhI�y}fja� G��a_@��^��Q�����M����E&}R��T��7�,L�pS����l�c}r+u�r�{�{�]�5������(.�&�ޯ�	�M`<f����A���Z����~{c�������	"'ᬳ}���67���L��g��ɋ�ɩ���%��Q֝�&;/��eb�m͎���ެ�WZ�5��?�7���|y����HFF ���>�Nm7μ�a�`z|GB�J��v��7�$3-�i�����m�4!�2��\�O��x� Aq�J�m��$ͻ"��+��f|'�u�
�6QH#j�r�QM>jV�m� �<f�b�w~.e�ёލ �j��*�5-.g�1��ss\:�3�+O�|����!L��K?�m��
��毉��׮1�q4_/�1
	�&���yN�,�%C�F#/b��;�b�`��X����I���֣���0SK�b6�p��a��0�8�/����w~��wL�y��5�Rgo��^^�(ѹ���:��I�[@��Ո�a�[�I�ZӨ������j*�|/��x�\�+׺^O�雏'���dф��ao�^� ��T۽%��An�������oS]�el���}����~9�s�f����!�F5t|x�RI��L�F��O%c(`��A�O��|:\ɸH���7�&�X�z5�R�di�$��>�6j�������s��A�$ه�J�{������1�<�N���O��2�J��Z�6u��񱝟׉�OA9��Z�����|��lط3S�(��ӲK�NMem�ƅG ���=�jX|�URr�r8�"�&K��\oU���XU�O!���u��(~p�PH�|V���T�s�ƚ?>����A�)w#����nԭ5����LW���z0�0�"�8{X!~35�����~"%��ӕZbU��.��3���eKC�Ro��/s�i��zA��j�]?�Z�� %eX&�b�
�֗�����8�6l��J��� %��R31a��֞�N���IT`��]��Ĭ�H��W�j�2�V���n�h+�.���7)�ғ!�3���4AT����&.�7��9����~�װ�Y��ʢ���ќ�Ƥ�B�,ee��@lWHj��mE�	��G��3�.���\��EG�'�w�o9-�0��s��{Z[��C�jh�w���K����S�>��an���3��o�o� �fW�^�	��d�V����R���<��P�C'S�߇B�lBV�p�� �:֗���V%or���mݥ9�]�h�y��2�G]qndBs��L�FO�p�G"*���5ǝ����M-��W�|S������\�'�u�BQ���t��8���pu���˽&S����q&5�v�����Y�]�'��Є�w�ʒ��l�L�Ge�S�����m ���[$�K1��X�Vu�ϖ�Q2�R�g�F�ކC�ّ���_> x�Y�p��ͽO����ș_���fLUhfH;V#I��[1�(���IM��˽��B���*��C����߄z�� 4D�葳���q��]G����z�;�'���.ݼ���ⰰ�HT ,M���`����O�f�V�寍h�6^A����(���t+2h�b
�"����_�!�h�JYx��W�ϵNyo�C�nu��>B,ۤ6,~;t`?���]����M@M]P���"x��ۯʏ�� t���T�o�P���3�����掟��0�1���tK�[�۶�Yr��D�~-B�&�T�%�u�k����l���IO�VA��6T��:H��	�?l�$x+Ov���e�S����g.Mt�3��K`ͥ��J�/�4�N��}0�{S��n�/��YR����� ��^���@��7y'��Q�T!��o���HU���3}A��d���y��K&�l�/��s�������5w@�[i���~�A��� ��,�3݄���	�6�f�M��ק�X<��m���~�~��X0J�{3�D�|� t��H�������)e����P��H?��O�$���g�>��o�oa��s���I���h��#��|��v�)1�,������;c~�Yj��}b�N���vK3��0�O[?��l,�v�T�|�sy�x���G"7�5)X�O��jf*W�y���ﭫ�.������t�Aliҭ+�&j)��1NB��((��=q=��nR�ɦI���2�rȲ��j&����I߸2gc	���������H�y4bY9�����(��w�˾�t��j���;�k�`dx+���{M�JT�������Z�l�t���|��t��\��&��}�i,w3]�c+��?l%���m�b���9g?%Yv������LV�Z�HϬ�^	d��������j�J��k��x]�E�n�X�E&6c������DRZ�i�B��S5���ug��Z��'h�NN�0����4$����\.�{ށb�i���h��
�Y�2��Wr6뎥$��M�0�7"Z��Rs4� ��Z���O�88%�ʫ:�����4� �g�g#-��ڎrӳܾn�Bax�iȷ����`H���ϓ��b��׷�7�J"+/0�O���N���AQ5j-�ž4��y��xQ	���$)��.�?�b<�2$�>a[g�s�����_��:���zZ+�8��g~k+�X!�*�_;��\������	�B/ �&��ө"���ZۂGנk�0��ڦ�_�KSM�`�>�n\�A$�mH��.�ؗO�C#.�AQ��Y��ZX��ug�<[;�ʴ+�?�Ow�x�O��VaH��u���⽈8 [觙�&F\JO��-�I��TӔ�[���E*�z��C @�	3K�>
�g��;AA�����\/�eԶt���F ���PmO�;�?�e�9A���o�ݣ��'rw�(�bA�֨<���Ű��	T���Tշ�sv"�x�UE��t�=�f\?N���KJ`�2�,5?���9������e)�7���P]�z��S���TAe{���>�{[�NYi��^�;8��D&��!���K���X�p_)����^��U|B��P�8�4��HڄT$��^�)<a]!A�7�QC6�������M�f���t�O	ib<�����?�6U���KѸ�t�k���`�%1+E3�`+1��+�d��xu���}��j���$�L��
lwH��IH�������5�=aݻYH�W� U���;�ꆾ�PE>%�*�hV��"L��L�K�!���3�}�C_��7]P�L�E����D4<+�Q��0�^yX�Un/��e@y͟o�B��V@���k�6�t��c�4�S�_� �!���(V�<��Mhh<s�!�t����$��6�L�¬34��$���!�'P�D��nm�Y�|׎h>��9��ƣ�Q	���5l�^͝˝n����*���M��s�y�Ț�<��JA���zKP"M�Mm���z�7��8�tA),@'S%ѕ��,*f�����^�����Xz�2�P�DT����.7(����e!X��ā����h��&S�����@m��Ra`����G4��	X�����썶p��[��ZQ�0�^G�l�E�����Xi6���Ե��a�"A�t!?���y���C�M��T2�]�6��"z��9�	xA��F��lq �Xx��X��2l�c�Hkƣ����5��3���.�J4��u�Z�����i�����]���e�`�*���A)/�@B;���H��9���9�L+�o�T�����B�f�^~W�I��M2��CZ�L� �U��E���dqM�&4	Ln=W`̮>/[鿜��2uqHQX��=����'�3����#WV���p��Q.���0�c����f�L׆�)ɗ�qv�70-ND����?_���oc�������+�D�5��'����V/��=�ً8��xy�=	ĿY�4S��Iω�ױ[�?��BY7�-�~6��n�lyv�Bc�pȹ�S�W=����t2	����hQ�0�S0�[U$�\���V+����Ի1�`��/�,y�y��,�.}b�ߴ��6e�@����%ˌ\n���,�~��a9ޙ]Ow�!�l1jN'}F6%ڿ�6�M��/��XU����Q��ʸ��\�8r�z݆�?Ӓ��R��k��3R�h>��'�N'�~26P���d�5�t���nL�uj�$g�q����0����E��]LȰjF�X��_dB�����K�w0�Q�(���/�m��y�uQ��V���M��Ѡ`-�1̏��/:��"c1n!K8�I��*�	5U�����l�L��w��x�u�Ug��v���VZQ]\'DgK�]���$�T܏��Zfh��U·�L�E���\����M,-�HӡtǱ��2c3O>�*5}t�SL0��'<s�hB���>H����%ѷ(�H�V�7l}n��XE<����~mx�n!�&��Nc��7����s�b]#_��m`���J�����(�{K�����6p�F����zv�������a������t�l�9�ǍͤUԺB�d��U��G@�s�h�6�����4� y��H��6��Iȓ}��ލMN�95��Qұ,\�]���fY�yA�������zB�I�b&v]k�=5�[�#,�^�(=IjjSd6��:�b�^S�RR����D	�~|��l�* ��!pB��h��9��A�ԗ���E{S��E�Y.lZj�H��-o;�8J� )��gL��$�8���D� ���X��o�?�?�����XL9�����'���Ŷ�S�5i��Ki?�b�ZʑV�Ϣ|�t�4N�<��z�|G�����'ex]&�V��C��#�t���;W1�a��֎�ݝg�/6�[O���}/�_�<
.�1�җ���H)P����i��-��t��Uf���t���.��9t�J������`8)X�i��F�џ����Ki��{�P<��o��@E�' B�H�k�|�?Fp�B�a!���鏟�1ǆ�{O����\�~��K��=E��B�AǑ��]Æ�=u9K��Ǵ�x�3�?y�3(�4�,��B��!H����H�I1�I����r���L��ڙh@��9�	�g�A!:ӱ�]E���"�����)FeTdZ`����d���xR:�\��me2��g�h/���^%�A�Vpu�"o���䉈�][4����X�l��ѕ7��qG�T�zd�$��|4="�wR6K��T.�c���&;�Y��xb��&*����ĸ��1:g>_O��K����?pg������'��:���x	�{���z��Ͻ䃎J,��\Ř�ңp�UL(v���j���7���$;[�/w1/�A3�lQx��������`%�<�/ey��C��_�� ���]r{�!ou���bM�%�Fx+�+��8�K�3�ML��S������h���c��?Ѭ�:�[�7�s�P��Bw�a�I���g������>c籋(tl��W��x�5�^��M����r2�Wm/ @�EU�-1��܂�r�ՐM}�v}9l�iB�P�1_^�ȥ�j�Z��+8�5�kW�5f���!����l�վ�ǃwZwY�eB���GH�%���A�#�<X�s~Os�s�E�Hf�!cL����l_8���
���ƒ.T�p̶����͹��UN�}�gߚy�&���%�F����Ұ^�Q@7̸�����u�X�Y����Ũ�y�T_�(R�TD���)u��t�!���	v�9��HZ\e����c[��>����uq��|(��iO!�R���8%�	[^���C�B&H��H/T��&[�/��Gmk�s��w}�N:�c����� �fIrZ͟�X��S�˫x��Fep��'�� ��r$�#��H���Lt�MI����r�ػ�l	���bl昳\�y�.��s��%��a�젾!�s^/�J�V�ݜoZ'
�;o�{��a�!(�MN��I�;J�u�X*$S��#�/BF-��t���˂��cg̽4�y�d����9F��2[_�N�j����c�ź��' �k�EN+:���v b΃��ƞ��,��C��䧺���bR)����]:��DV�2��<j�3+�}��V�/���.�)NpW�����y��G�|��kևю^���jj����"���!y��h&N�T�A��aL����Д��E�M��k�Q�	�ma���ȷ<Hm7ٛ��Oܨ�R��w`��D�yF��מU��X�2ig,5B���Rۓ:e���3p�װ�y	�TFC�otJ���D(Cu������`��6Ԩ6��w~Ϧ���\W{�IT�|�5$\�֜�x����%�l����3n�9]�B�/�[�au�����G��W28ԝ:P��􀲿��dv=	(Q]ˆ�̥�|;#ЛG�t-hw����"�,��ؗ���Y�!��(�+�Y�O/T��Td�c�����V|M�*^�Z�OcJSNo~i�'>��;T��;�ؿ<BF��j�@��.�1,�������l۫��2��w)k�jٿ����Mg�7VOX�)_R�p�<q*��۽��K�������:v�댍>�%)s{��8R����א�
��R㫕�Ɲ,��.��!��t$yfI��y�)�ϧd����H5� y�/��"pN2�z�jF�D�^,���;�G��#�|Z/��q�Y���U����8"���ЩA_E�Vʄ0I��ʡ��V!����c�h^��������9"�1�NS���Rʤ�Fqُ�� �����b'[T�W�)��ʢ_� Ӏ#)щ<�:G7 '|�����&�T)�G(c��nZ|�����w���g�o��T�6�~X##�3�A"�ԣ����%�W4�/���E4Zwa3*�� �T$I@)}s?��_��h�/y�(HߍOq���6V4����r}`m)v���$�j����f,�z��؟�ǲ�XYm�y�est�oLdq��%����x�˿!�Ϗ�h��E��ͣ�B11�&Fء�i��O�%��]����R3�
	�<T{�k���ȭ)Y���%�l!]�-|W�"p�{�AL,~��_�s�\~4���e����{��m��-#v�!����Y�!��{�(��|��&�� W�U�I�nZ�� ����;�������~#i�Mϵi��bfl�-o�>K?)���$�n+��䅴������X	��L���A���nޙ��Ɓ�i��N�X�mk�X<���+��v�;b���4����S��>�����=0��I��@H?K�D��#,,���T�TSe��m�[e:`HX9��E�<�K�@ĭ⅋O�[�FJF�Yp_!I���E���i}d
���qd ��MSD4c��<	eT\*�
<��qC(�I�6��(�R8Ii<�S���w�|8Hi}
sA�CF�|ü��j����_��ܣ��A,��]�O��*gJ_������b@N�5��1d�e�+���M����1/!��f���O8h�)�G�N�n4Θ��.^�tVԬ��C�p�~�>�b��ewK��mL^��Eﳆ�~̺W7��o��j�?� o�F�q�^Q�P)G�=��X.��<� ^C94�5:)�*g�s ������ Kx�X�e0��XH��!e�j4�߶퀐�����Z�ttt]3JfSi�+���V/?��tq���	[&��.6��:��_��o'��->�3	E����N�e�ϫ�S;O��ܕ�ʰ�K�|5�b���P3��rGB_���W�&���o�r$�\!��]���kF�&&�%�'2`��5j�4���E���à���K/di3-N!�'�i�nRaf�;��/���;p��}�����^SU.�6���:v"�p-p��%�I�x\g��Q���G-�eb.�M�Y�'q,���wj�Nb�9il���W����8�1�G�V��].�_��mSs���h~$��+����BS� ����٣���u��uY����@ $j�N����R� �c�\�ϙA3r�/Bv���(��p�d.~���l�Hd���*�?��l<\���?��:4�k��'�[�t
N�����!k�9�`��Bԋ�E�NZS��Z��
�Q��0ey��]�n�UQC]I��~�Y�:���Z�e+���G�z{��BA���x�%a-�����7�,�-{�����>�Sс����@.OQ���"�ߪ��GL�V��Q.X�6,H�E1:�,��?�]��n̔�R�SP �H%vˆ6��eF^����=��W�m��*{#�I�Xb��>�|ĭ����wa����ED�ȫu[\����*G�Gv%*mkΕ���O��z[9���h���tFHy]U�=#ַ�Zg���mVW2�A��Bر4�)��W�tUH =�:vGySd�d�8*� �bb;��;��]���!�6þN�m�D��U���T>�ƃu�	魖�.H)nF��)_�x6���3�
�ztu��vq�(�΅�Y��^Uf�g���o��L����5�����
�{6Y@0��WKc'�sE{�%�s�������� :d�]���P[ύ��\�R�M��-�Y�2	y�/u���D�Q�hW������_�J���bF{�]���>'\��5`���&9)Z�f:�?a����������5C��D��A`2��&������R+qki���/j	�b-��/R�\1�O��m1:����'\YH�>ݑH���͸x�K%��ȴN���pI�khW�Ib�O��"̺�E�_��kG�k�%�����Ô��b�Cz���1J�:z��3N�h��w�{��N.�̮��>%6���(�k��p�HK����ƜgR��gZ�x�)����(�fy��/������T,���e�Nm�|p�v��9Gz���DW;�T΃.R��	feNp�2��N�Mt��\�"���[�����X�"M���Z�BZD�pe�sm �"}�j]6���|�IJ8�:/��t2�ϝ@Ԁ���6�p��@��G[@x�b��FEO�����lo��ϒ(���ۖ�ޡ��զ�ºoNcޓSS���WW����wȧ���Q�F�����⨲���7�����̽꽗E|�bbyxsH��wZ��J���̐�(�O�ͼ����`��]�en#f'J[.v�l���XZ�4:u{Td�8%����ɪ-�-~������]�dLo���2�D���/�B�����E_c4n}b_�=�����,��mw�!�����D=Tob��kj�-�|�>�>j�c��M�d���^r7��b<K<�$���N�p>��3�|�6#� b՜��yጘ��oj��pu���'�DmP�)�<�|i_V<K� C��M�����-F75��3[AC7�%����L=��p��1~��s.4�۴��2��~�'�Jw�$���S��.��E���W�NJE�1L�=��l�x('j�FD�w2d�����`�]\�9��bAg�*z{.���JA�Y�%v�mk��-�w��J�ۚ4Ka�
��y�7���z��[��R_$�s�T]�.1�{��kKZ���{cq�r<�KC���(�.����A�F�`ơ`Q`�7�A�z�+g����H}Q�G��* t����6�R1��(8�~d��������@�@�$���B��q?��7Ñ+{#}�s��+� ��И/�7���������/8q��=Ƃp��u|�.�i����.���#��Z�f�9�@E>ȗ9Z��;W��	
�&Qx]@��΄���<�]�!��,X+{҃(eS+�l~?�y�1�rGEW݆^�??�@cLLP�0$"ҷ�?nrDML��H��e.�A���W!�%�	k������Oc	�x�B�u6���3��k��f�m~�[��'�9�",�x,�����v�q�.-��g�_�c��~��k�"��g�l�}�a����Nqh�x�g4Й@����v+�p���q2VJ����y�<�~�3��ѫ�pM+w�p�B��_^��Ā)WK����MI��I�>�"��⅛���׵$P�>�4*Bc���nL�̎�t�F3�6*@(��C���� ���䍞�|��7Ѳ�1ZԂ�[�_�B8�I%j��*�&���P?YT\��e�L�u�Ϫ��7+P|"�Y���W�v���zx+]�W)�h[�1��ܕ"�����(=��L%����y�ɀA]�OM8�	%q��b2�i)��
����8R���m�V�@=��z�:b��=�s����@lY�
�TR��<�K�`�����`�h6�]�	|Y��|�0�?�V��!
��$n��n{��P���4�㌐X4��R�o�*}WLT�>[�����ۤ����%5 �21�v7�;Y�k�f��@`�J�9�d�Ǆ.��|x����s�7�Z	J�t=fV��5b�;��(Fn��v�;g�@��0qݤ��Bd��;�M����|�c�O��֑� U�@�\,V�d��������A6�z��Q|�ڪN�(9�f�Im�Nk�j7�X�g��M����B�
��ڠ�"�7b��:��J�AB�{�=���ǉ�ݵq����c�$V/��J�pŇL�琖o���$C��s.
�ۨҩo6@�4����sY�Y�2�笭������.w�)��ꍦ@Jl�ݮT�M���ݣ�n��	b�p����t�nt���>��R���.n�U�� �l7�A��a�`I>Č�˻Cέ�2�n@�o�H
���|��Lk)�8Κ��"��}Mڬٵy�1�~�S7��{���\���w��������,4NM�_qm��^>_�U�Z�Y�X��l��~�d��tL_�iUW��w��U`9F�6�����qݨ�BaG��ғ��d�u�3�C����P�6��J�k j����ȓ�kg�����8,�Rx;� BG�������R���B�hm�nE| /���.��SSSN=$��_�b߹w�
~Y)�M�B�κ��ܨ��?/�O�S�s�oZ��AO���W�^#ܒU��3��:������G�fUQ�M\��,I�������-y���%���?�N-Tnj��7+7�T�7�\�v"d�ʊ
1f��v��uS,f��2�o�.;��͠`0L]2���+3����.�B����L��J>i,�U�����/dKA-�v�����B�I��
�1<�^S~��N��=�/à�#��N����O�\����Ь ��xb�܂�٥xP�{V������I��������SZI�g+n��1϶
kҠ�)q֙�]�p4��-Wf�o}ī!��WEs��֌sLE���L���2A�FD�ٿQ�O45���^�Q�L��i9� \Baޤ8uW��L�s�d��qNUS6�JiTgT�ܓ"sa-XTOˠj�L�@l1�VH��	)�W�ΦD۔�/�lu�U���i��"4���SB2})`y�Hl���Bc^V�<�cpJݩ�`���}� c��c˚��7�S�BI��"NU�G�\�VQ�E+��C��D�e%�qz	�^;[v�3��I�L�C�q�YHf��rQj�`���z?,���T$&�M^{���n����s���E���B�]e]��/��}i��\��[\����*kE���B�mcG>��D\.s�H�����P����u��q�mAܵ���)q����-պ�M�����q���TP�;���ʝ�;~���)1��)�%������3o�֐m��}����#wO�L��� �vT�~���		��? ���l'7�W��2 9f� �4[b�z���)%ԣ�{I)����� �@]��#������!�-���J��c�+�%:�m��f�(ez�ߜc�YвV+>���s�u�fn������I���Ul�P�)�ǋW��賰_�2L)ʵ��Q6�Ax���gw�	/���M���C�ݓz�L�S�'�x\r����×f�9�a �Q������FC"A�N�b{�=��M��`�_*�eD�[J�S��Ԁ�Vdg��9) �EG�C�ފ	w��eAF�a�I��!��� k��35c������D�k8՗	R��;�.��b�ڊ+rrl�Р�
	8?��g����x�@�)Bl�S�N8!�?Lѕ�0C�Ĺ>�KN<����x| �� �+^������g���6�M�Y��0Q�����we�Z�@�0�
�yӛޔ�w���纍���u��s�'�9�~���W�����`�����1xŊ<��L��9�Z�^~�Eu���r��}��Ҽ]O�/���ݕz�V�wݞC����Q�kH�@먭�FO+�� �#������/~q�n��D��Q�
XVҳo�]��Z]�r�E= zjq��1��@N+c�� `F�S�=u���q9��Zt�����O�Ld*uۉs%^�v��d���Tb�Mh�Ü�!q��Q ��m�C��0$Y�\88����~zf�_|q>�{�J����ʤ�Y& C?D&|��_����Ȁ� �q��B��b� k�<Ϣ�Qv: �C����_�>K�<����`�1�'�@�K�ӷD]�<�(�L�����!v�$ �Fθ%R��aׁ0Lx����h��=5�gR�#*=ݩ�ڗ�w[c�*��2r1mrT� ܞ�KePpב�ȱ��S#6#��T�
fZO�0�3U��t�i*���L	�Q*�ؐ�T��
�#3U�3�2��Vj�v�H;Lq��Id7|����wU��{�Ȅ�n�^�|�3�fˆ�@��9�����$�=Lլ�� ��3����͟�ɟd��������h7���p�'?��p L������
�I��rl���r��Z~ٯDCv\�HƫK�2+�`�H��"F�dR4���Mg��9ޕq|���s�,77���'<;�Bݩ��|ڴZ�.�#��~��[7ϫ��ݖ��&s[ޏ�]�)I�49NOdU�21�����kF[��h�TH%`d :�"L�LQ��Y�:���0�9��t<^GpSs�7�8E��c]�n�Yb�f�L�>��U9Ǻ�םj�Z�2�O��3�,��M ��h!.���`��:�b�s��p�3����&�L�Q�����.���Mٜ�s> eyZ�O$��K� E�J6:�@���;R�%��Y�83^)��Z:�xvC������F����\���rD; �9G6ie�����t�v�:0S%�6�{��QV���e���eW�C{b���vU���d:Ʈ.S��og:��:y\��V��} 2��ѣde�X�W�.d��	q;˽L��i��_@f��l<�3��,��9ޫl��g����8������Єa�0�hw6gu���~�j�e��z���-�	�@�=���.�&6�@]M�c��ϻ�p�C��e����jh�:�D��||+�����j�[��s��Ϧ�(�	�o���|*m�
ǲ4�5<���'\�����#9R*3ǃ�d�ѡ�wesmw}q�pDs�����ɮ��+����eH"�>��@x�W�Y�欎�������m7]�J�`ٲ�/?p4��4V�9 ���ifG�*owꠑ��iL+�a<m�	��ɴ��9����R�w�39��X���Fd����9��3�@����+��e�Ɠ�{v�Fv����b-����J���m��I9n,���~�}Fg,W�]����I�^$�)^�N/PD�HA�qz'���1����=��bW�^f��ٛiVciP�-_��h���>���y噒}(Cd��i[ATPҾs�/�jH��r�w�R�Rc9d����}#�R&%>�,6J;��V��?��q��LR��Y����O�]���p�#�n�|�p^���1'Ǉ��3�&G��:T՝V��S�q	�g����f�i�H�S��2�3�g��_�~��h�ZM�:y�v�S>��?���.�I�2�`�{3p�vY�q���t^�R��ؗ���<I��x	 �|Wէl<�|,K`��͑��s���f�`�mF0zw�R�̺u�N?��#o�H}��ʲF�	�� �մ��E��)�^RW���E��hd��v��Y�x�*�����r�:�SnU�~ou�V�G0j����X���#j�婴���-@Ff��;2j���Z�M��yO��+���X�0������3<�(�,ʤ�2�7��U�� (�-�c��s��n�|�p��ㅨ��2>��SfZ��y+�G�h�܋�1LE)BQ>j]�u�V�G���j��"�+�ɛx�`��f�
|Zw�f�<������FS����Rw*l��L���7��T�]�����D@x�:δ���f�QS��E�7c��]��}z���-���c�N�X����""A���N�v`�ʲ�x���׬YsZG��	/������/oo��;;��c��Z��<FR��]5`����`#����>d&��d!w���ޛ�Kz�����=�<d&$@�à>8]8W88!��H!�	(I��4�� �E�0	����9W�<xQ<�	��t����I{���ߪ��~�vU��ݝ&���~�v�7�o�w�����w����C������Nސ�{��4�?���u��Vq2Ĕ�|6i�B@��^����`x�&.;��>y/jy>c|v�t8�s�i�u�F(�Lޙ�Z-�z��R��J�Z�>z9���8.u��aWX��b��vw�*��6\)�B��w4h����� ����;A��ױ�;󌶣��+l?PF��ڽ�a[)+,�x��ږ7��E[�X��$>�P�U��;N���p0�r8�AaP�;��fo�?�~%��ˤG��L��a�e��!�JNpƮ�jc��_q�[�V�;kl��OW4f�&wD�I�v��A��{��M#�+<�Dt����r�2��xm��GOS�WG��6e1�[�v���	n�;��C����QX�������̵��8ײ���SO�N;�����9�t�DHT#��6��T��z����2�;�t�q�{sv7IPt�YZ��M؝��
2�����בN���j�2��x~l_;{���t�lo��{rڹ׋$"��*��vsH�bt���k��*�����Η, ��6]�f��ދ���G�T�h�����L�jc�����O���\����0{̭���?]�i��ARw��lg�n�j��޿�`��X5gn1CЬT��Y�u1�/�h�Le��.��iԢ"�Q>¸K+լJ����^�J+ѐ��k���wΑ��y� [��,��St)�n&�<qW�����ò�Z�m�W���w��q��2��`�إV3�F��|��<��z���w��P�o׎V;�z�Z���c���!��\/���{Q>�8�]��22m)��=��k,�m�Q)��k^[6(��l��`�,��F#񐱎���^�l�2�Qqb>�a���MY�{�s*�r�HHr�V��r�V�]w�UW�jI�����;n�̺R���Ä+�RzԣN�L���l��/N�H�#h��ei�y!8V���e�s��;BEG�!�d�ܨх�]D���&�.2i��\)�1�G�^�@X#��x}^܁,v>�5���#덁�����An�K��ۭ�y!�]/v�R�ee8?��^b;R'�(Ld��@��<Z,�'QI���c��K��!���ǳ �<ܯA OY��m㦗`��b<��B��s�$>�ed���G�х��R/r�~�oJB��ȑ)K�|^��B@z�AY�s��&c7��"P���|�dL�RO���Au�wl;S,�f�v��M���tZ�Z����v�EK�O|�N*m����q���\5=�'-_�2��-K�{�/��ǬLS�>���rG�0��Ep�x*������������.�hV&�����'S�Qʘ�a!4j�S��m�N��`#;���\��+�� l|�7x�r���y8G�F!����������EcLf�r��B d��c,ovfoԜ�VK�@-���mJ�F�tZ�Vj�j���p)M�v�n�<Q��R��g��ZKs�-&�Ʋ��q��Z8�>�ff�a�A�}�iD�����Bo�kE��s��%
Μ���
��[�Bd��3�+�[��a�ڼ�5�=)r�������zQ^��Pzp�n�Ȁ��00�%c�a7q��wq��{S�uAuKH�	q�l��v�Z�^��˖���8���K��u�KW������M˦V�5����^v^Zw���h�S�Ioy�1��L����l��	����IK47��7�^a� �ph��Բ��z��YfJ���Iৡ�%�G`���q�?��@б�.��>sv$��q� &�|@'Sj�H�����{$\���`��9���2�����K=��d�m���s�Lw�;��� ��	˝Tj�ScvO�4gR�4�j�N�R
L�?��� �K�T�J��e��)�jm�9m���|���Ԛ=�;�8;��@؝ǩG���DFL�b#�=�.��Z8�>�od@Sk�ހ�KP���~a�7����=�D� �;!G�9'�+j�(qu�m�p���ƿ��N23�گ�Z|�%���ʖ�CdO#�}�g��.qv;4�&�-�)i���C�R/�P���duR(�,�[R���sL��ˎ�o��S�{V��I�Ӻek��g�����J�l�9�l��
uD�*�
#����/�A��R1��#}�@�zq*�J�0HbM�9ݱ���0�0�s](#�I!H�����8g�w �IƉ:F��4�ܫ40�IM��Y2���:-�b��#��?FFbor7ctb��Ip���:w ѭ��)�k_��\>@��_�j.����G?C���g���x�X{ww��>�y�/��?.�����4���T�{_�vfS���Cw�T�ו��y�;�SO�e+Ҋuǥ�D-�|`w��W����1u=將����B;#O0���P�7o�^ �F]GF��ɹ��ljp�%���A�w !�ƽ��9�k�17d�K��#�a����e�l���	�-����}�k�@�?�����v��v�n:� y�k�naͤ�$g��@���7�Ŀ��/���u�s6Q8��s���ɓz����IEo��@��D��z{^d�⊍K�;�W]s\���t�=w�]۽s�Բ�43=��_{lz�K_�V�_���_�����D`o��N���@T���i���A�L�l�� [#_(�4�����Ї>��R�1cr�4�>�bg�,��Ʀ�0�j�AS��h?��?�wQ?$����<�0eư1@� &�8�@y ;�b||ϳ��]�ʝ1�5��n�������
x�	s`0�3���9i��N>�Բ�bq���-w(�g���Z�6U:�Ԝە��ܞ�voK��L�4S��wC�dT�Bڪ�Ruٚ����R�0��d�g����O~*�y`W�*2�4Y��obx��{k��`C�Y�\u�U���漋/���+z��&��n5m�?ڿǩ�9~W��N�y��6b ���������}�O�ց^!yzق�~*a�8��>�M��A�z����&������ۋ.�(��+��r>G��ӟ�}0��乭�a�T$_`�7���_n�Z�J�z���.wē6}��t�Mo^��g�n��2�RJ��~��t��ek'�?��?�;��Uw7j���ac&>ӹeY���\v� �mDu%�*�
�qC�#{>9":s��rC��h������p�0W\qE�����2'TР.���h����y?L���2���svW�%�<���tf�x���)����n�|��~���;5�~9p.4P��戈Nw���=3�3�} �ukW�jj�NcWz`�m����4Q��r{&����F�of~�rjWji�]MS�O�ם�Z��4ۮ�=Ӎt��@15�-1?�K��s�zPF�3	�ِ�v�=ٰ�}9��/�D�p�����'�5��0a�Jr��y�X����c�3F!p,&�7  �����D�6��3S.�4�ͩ��:����U^�n�����DٰU��5�\��i-���og��>���c�9����{�2�mL���� "ЋqǲpH#������2����\�iӦ��l�r�;�5۷���]_�K���w��?��w�ȳ�j#�QL���]-K��ŀ޳[* ��>8����7\$a��ѝT�<�Q�A��pܓ�`��@�k;� �E�t��(����.L�Q���t[-#�lE�ar��<��S~�2[�Ȅ�;����� � �lي4���W{�9g��kV�j��R}O�ǖ�س#MTfS��Y�n��@�E�Ze"��Ժ����N�ʊT��Ү���k?��y�� <37}X��y�`�.v�� a��QA����:�������b�N�	���{���\_�� ��7lؐI�2����� �eP@���r?���9���F-�S׀0�� I�B���b�S��(G?�����_y��z����#���1�K��u���;���hh��w�<�v��n�Q/������a I��z�D	ڕ#d�����O{��r�Q��S\��q ���(r�$�����1�"x9����սa�L��U]�a�}d�N6Poh�	:. Lgְ���k�M��e���.�4N�c� a��{Lx:��Yg>��{���r=U�3��Zy�-�$=f�e�<�f��ij�Ҳ�'�fuEy���    IDATjt���F�����;YK��Ls���ʏ��Ud�9����l)�0��Z���u��g��Äq�e�Ev���XU\G&s� �er�~�oܸ1�=y  �F��"���[^���~�ٸN�]���ס��s�6H�ֻ�޹�[����/2a۪�^O*�%c�yb���/]�}�KW���(G��Z�利5I&��G��x*]ȇ�� !t�8�{��g&,
tL��^���Jd�g� qɘ����?������KV��԰�);F9"2�x\����p ��f�6�=1^��	+G �c(�x�;�^O/�[��%�޶�0�VN�yu\^��`��3^�"���J��g���Ք��� �J�SOӭZ�\��4�^��Jiz�����S���v���j�?�m��� a�� �@8�罅N'�,�r0a^xA��7Оq��Q�X�r����BL8�����R�0����~{lSc�x���{�gF�H�����C�0���w���c�0��@��@x �B�:����K������ߗ��q!j��FG�h�DG4��R��b����3�<8��m�*��|����W������?��yGe��ʥ����p�x�2]EA�@@��	;"jx���"ƀ1@ga�(����a��Z9B&� g�#�ZV�a��.1&@8�NV�#�h�y�E�1=���rskV�j��R}Oڵ}Kj��@�5�Քʬ��p^�����J��=:5*+�\�H{�&|mᩱZJ�V�m�Lx���G;*���d���+�� ��V,[�`� ��0a����=�����*`L��Ӡ_�=��<[��1��g w�8�#���b	���w�0�G���g/{�U�~����9"t����w�ؖ[ߴn�֗���3��!G81�z��Q�T��dD��3q|<n�F�h;�c-ch	L�0�^A��R�V!��� LF��C�T�`b� ����
�v��d"�	kP��Y��݄	�LN��	+-��9�L��}r��4��)�w@���v=�K	
L�e�Tji�UK����?�µ�go�����/�tA���$���~X�/��E9"�	c�Q���)DQ��Z�N���	s���Q�9By��F�҄#����
��Ș`c>��h��-�&x�2?䜋a��r&}����Z�HȜq>K�;D���> �D�r�R�0P\)W>�q��Y2&�o�r��mY>��	+G�	�<����y�Atw�Q�o*
ed�a�0a�)uc~G��	#�S��-��&���l�P1hX/S;��&L��LX��r� ,�	�	�|E�ӯ�<� l]'�# ��R� ̵��N�9p�/f����l��gow��61��# �j���s��m����&<�A�&	O���=}�SKӭj�:�4��ѩQ]���X�=3�>�'�H�wޗ&�*Y
�kD�]�y8�� ��'抚0Lx!�s�	S�h�21�u��"fg����BrD$&��RL̙��? �L ���!!�� �=�	�Y&�g ��N���	D ۧ�=��Ȅa�BB��	wCtK)]�eo���x�8�kA
�_6]��v獗��~��k:��r�!j�	3� �0#��ZL� &���}o>o� ��R����f�a�R�Q�U2�Sa$�\ef��n4A���@g6�� �L�Ɖ��QR�����K�;1�=r�W���R��+>w��$%���e���_si_�/�gz&�zr�Yg�t�Ks�i�@��4^n�rk�|��	ۃ7Y� J�SK��JZ���4���ԮN�F��=����O\�vݿ3M�Є�~�8���]>+�	AXa��1���A�w���0�	h�Z�����W�l����8A/�&l�@(�/@� P�/�cC}�����%��`BX�K ��=��RF��sW�ƍxi��s�� a	~���.��%�n�d��7�}�D��Fs.k�G�X�k����w�9/֨כ$���>��E�;l���S:-yT8�'0�όV�D�<u����9Y�a@
��B Lc����]Ӹ����;\��o�9���c�+j�>����\ <#*�3�%��;�񎮜#t,+��,̆�}��O��O������"7�w�m}h��c��@0~<
���Q��� ��^���k�涛k�s�=���H�֯J�V+��{S��>�:�T���$=dI놪�"�Zf��jj��Ӳ��R�6����|`W�����������R�3.�E���6�J4�Ձ�� �ع瞛m���f}��`�=�~�d9̫@����*^��+%$J}q��r��r��/��x��!MG��^q�_��aꎸ}"���g��7�pU&�|@�Uϕlp���:+�5}vA}��_�܉I�&�ўMF_a�"��[��Vf�JLeT�奍��L��/a�s�  ��+קs�9{�����F��P4����T��K�g*�����6�����??�Ӏ�Z��!`иѭx�k�PG�<*�5T�����p���x��v��m�c��ѹ��+���3�����q�����3p�7#��z�wup�� v:	uI�v"�r�,�@�R�B6F@0�7��l厲wzw*wHu�L%�O�	JC���vzrn;uJ�t��.�)͗�?$�I�����gg�\�,'�!qζF����开ðW%7�L��Ja�Gam���{�mhk��[��`�\��z\�T�s�|��U��|����+Qh��Sڟsjȁs<��(a�+'�B���;/ u����_�k�\�?$��B&���	��sR2aޕ4)'�f����	� ����m��ǰ�{�	�G߻�es{s�	�	Q�'W��swo�'��< F�ȃ�E�Ӈ���z��X5B>�|�+�7C���Dy�T@9�YN�`�#�tw E����BY�{;���n���\~^4�c��5*#8�g��c�%ǚ��e�<��kG�<���,Nf������ێ欲J��;���r$L5�X�2Bml,��͜f2wn7G�3(3���R�CFo��vE�[#3[9uJݝ���rg�Tx^K��l6�� ����9��;_!�[��ڹgjF}�,g؏	��I�eb(	H��r�e���1#Iq�s햿%�c��R
�k�>��@�}�Q��s,�IP���2ǵMٵ�9��dE�"y�
���s� �sAl�ޭ�'l�믧�a���.�b�'\��u�-7_�n��,�OS��e*9���5��;�� L��
$8ډ�ج�4L-�M������H�{�~��,��Ÿ�[2p�<�09�k��w��ϡF仃�#�����������Ռ�P4b�se@�!2x�`Y)�@�=ޭ;����*j}�2c�Q����dڳg:w�����]�_��J�(l�����xNi鋏� 2���r7��lf<�̴�e��i�T��;k�ژ:q�|�w޵m����i[��AS�4�^+�B��-pm�%@�o%��mS����$]}'�<���8a>,�K�����9DGy c0c�/����"������[W^.��PO��sb��˲�񪫮���SNY���·�t��w���>}4 ܨ�Ҫ��U�ze�#����Dt ����o�v�cX�#G@�u�u�96f���e��m�y���hn��Q@ΑLY��y���)�=���4���"��Y3�]�0��s�G��2;hɠbB"�*0+KP&Yב	��b�֭�
p��1��m�x�,GĐ�ٺl�,h������>l�=�z�}25�����fNٓY��a�|􈔥�;�M�eE�q��H$M=M�\���i/�BU��{��s�;��2_�U�e��-Cq@�?���j>�y�s�9'�>Z,Rk� n����\�} ��O��&L}�f����,��d���F�	��c{u��+����3�8c�bLr������fn6�9N��/H��N���{`>D�Q0����o�[��u���+�뢱2�����?�gBۘ���'?9?)%��9%��&	���$`iL\�g�E���02Y��׭�ÌP�Qɂ��80(?Ȗ�`�r>��f"�y�^2�AL*{�;�ZwϹf���c��ɚ-�h���p� A&��[���;ώϦ�e,ԩw�F3U�D�/�AD�0�M5��Ko� -KS?��M��ڢ����� !����%l��%)1.��t۲ľ�v'�U��k��/���,- E�s=�(̗�)&�ɦ��+�����,�L�9��6�tؗ$�(��L�{�b�6�1�ܰa����~�]��<�>��n��<@xl�����E9�<�����֣̄͢��i�bG��#3f�W��ys`\(��a� /�1Ǣ;�-S�0a C��VrԈ���s-�@wD�����Fg��*���!���6��;��\��VR(x���a��L����>+�*���@�� �����x^|��k���|4��֟ݎ��N��8���gV��:�%2�l���}麉���C�8�AX�l��HF���CQB�]e�\_�I[��;��l#�g4�'��{�����ne�[��]I\��,_L�ﵰ}u�P�c| &���|en��}�c h��|�#�޽��� w�'�-��IY�񊃟�籜��Ah�!��,j`���6m�t�i��v�};��B˄�m�㼩ٽG��*�	31��lot���y�幹�A�҅���ő#dt�?��2aN cbε߄��b�fA��1�&�*�@�gu�ڭap2z��	|�}d��!:�g�3�\�<JCq-�����!"���xΑ�����!$�l�=J9�݂z�ϝ'�z�1 �;�ZBjH=�!�,���Y~�)�~�VsS�a�u�N��+��h��}ɬd�F���H��.��&���Q��DgP��^Ji��z�����w�C��r`'j���g��{>��ًz���JH�>��d��k0Q�¨�<�9��!I�I��)r�zDB �Ω���[Ǒ�Y/Vγ�l��ԽK z}������Y�����^��_OG=j]�7�R9O�,�D��+��y����	��0q'��s����x�.�O�8�1�]�����OF�ae��N����j]�!�ݒ����Ч���9�#��=�%�3�D�����' J�	|�A��'+f���$	��`@l19�9�9���A�_mI,9��7H�׿���9�����7.=fb9��LL�q�?�*S���Lx��`�x�1b��{dc���Y9�	��^3�?�����+0tm�;�Ły�\��
��`���l�N����?�:���8�4��Xc"��D��`�C��8̤��_�vԉq�s>E�2HT��IO.��M�6]��r��w�ly}�(V5�	���W��g�˫�ƪ�AX�(6Ha'�tK��t�8b�����o��[���ԣ���[����} �V"�l�8���t������9�> ��~�<�w8���m8������E���?��qz�1p�	J�?"&8�����b=쨕+'z�b���w5��u���Qwo{٪��Q$[�	��hPմs��4>9�(&ܯAc��j�`�:	e$��ް�aF+yn���5�����}�0.����}�5Qx�R���y��r�����#��?N��	n�6�M��~���\'���W�XLTw1�I�-�V�W*���#�m7�q��-/[��G��g"��j���6wg>��n�[���̣>�䟫���1��� Ց|�{�a�H��s��j����`<�����|�����]]w�u�j`��������Z���A��z� ,�ᤠ��N"F�̶U���,q����	L~�zr�W6n���%�# ᱻn|��{�z9 L�V�� a��L{oγ2,Ns�0o���9���+��V�P7f�~?21w ��=7�n��*�v�;��v�wys���q�r������a��;�j�+#�\�m$��(��|̓B�x������L���x���	��[��֗?�)O!��ȯ��,���nٚN�hw��Y.�(�u3`��[�,�s<�ai>Le�����1C�z��O�3�ar�~����(�@W&�pO���y�AL���_Gd�Ca(��X������g���ԐP%�w����3���?��������֋9�@��SO�:�^��A���ׯ�~��W6�fb�ݖ����Sg��[�D'�%,6�ofTn�+��=��w���T������[̳<���P��@\�{~̝�x���=����l���{��#g>���R�[c��,=Vف>�*��t{@9���k�S�ʠ�)�r��7o���SN9��Ŵ�� l��r�ZjV��)�R݅X��������X���`�����KZMFjK(���[��:���P9b1��	ˈ��b�q��A���\l{ŕ'��+5e���D�$�i�{e��_tԁ�ㇳ5��`��A�\��W]u�yK�y�ܭ7�~��0��c� �q9ڒ��\��s�6� P+��$��A&2�f�{8�ȽnE � �� .�D�E���8Y�jN@��f��u�����)��7z�#	��M�9��;�a�Z���j�Ì��uy��/���F{;��v�#W?R�k@Y��t��#K!y�@Ў��
eCsK�7y]ȯ�>+�Ҍ�in�w��E�nQ4*W� �,q$c���0&���,.۞�(��>�F;r�!�m\F���6B�g$i(Iؗ`����0�o������谍>�p��(���9���(�H]=L��+f�1<�p�d(��G�ɑXd�Er/��! ,�XH��VJF&`��y!σL8I ~�0s�-Yt�#Ev��8�r��0� L���y����g�0,@�\d8r��8�5Pd��0L��~��v�1�v�>$�1��c�̎7l��VaE���U#$GT*��]y�/;�.VZ�ճř�@�`�	;��	�9+G�	��Ȥ���!�mGnv��� v��y�a�h����!Z�u�
�醝.�$� \.��f���K'��	o}q�?���F.�/c �����_�żݒ��ѥ��@8.m�G@xXm��P�@�s���� �0a��[��;�dA�/���~�����!?��s!D��k��D$���	Ah��u2�c�ڞ-�ɺ��6&H���5��r-�0'�L>�;������ƖE�^
͌k��刻����hd�<�Y����[���y7�
[���.�L`�bbr:>�Ƚ�ޛ�u��s}��VH���7�t��`�����{mٲ%��|��e[,⹑����q9�^�B�R�~u�,Wsq^\��O/-ڰ+DM@C�L�+������ص[w�)�p�B�MxII{p��?�Wd��X��.}��gQ�I�e۴;OOH�LܐN�ܾ0lb����b�PW�@������'��S��T�KʱI�a�&'|����`"2CGgwדN:)�b�c���W i\�]��b�<��>��d�@��k�f��ʕu�����Ή���!7�i�������H?��?���_�%�n�S����1���V7vV�Ϡ�f����|�K_ʠ��I��^���];{�3��@�\}��Y]�'��C0����֑�� ����]��^�i�������`��D�;�=Ԍ�e�
<ĸ�2[���g�gyt�W~�~!GY�C4��5�{�����ڇ�T1H.��}�W.]�G�!��H؋���җ�4���+ۨX�	&�C�@0�������{���
�H^�WdVH0�w��]9��k���N.����Q��,u�cZ'q���԰��ߣ���i�π�Fa���.|Da�,z�=��[-]t�E�q�{\�A��g?���c����3��_�u����s];����w `�^�'���9>�{P=Yp��r�D�@�h���҃���U����3�*��    IDAT�SG�`��8�/x���J��|����y�>s�"~�gӞ�lL)�q�^{mցy.�����y��;+��>�����g�4�m��詍b��# ��L��Hq?1ȗ��e�	c��: )c �aN��3t�p�]�I'g��a\�}�{_ޠ�� ���
p�U���5_d'�Q��X�����2b:��Yf�Y뉎{��f��D�'�k�젋����~^��^l�~��s��l����[7$m
�������K��F�SIF��͠�WN�j� 4H
�*���U�
S��?�4ݿ��X����yW���-�{CD(�r �F��`�\�m�b���p ����R~Ҧ��Mw~�����������?l�#��&�@���8&�KÌ�&Ʀ~��adweS��i��?~�{ߛ�p��T+���<kT�AF�q��s���b���xc��S�_�T����Ox�2����:0&�*r Mg��;���5�I�y�c���|�A�B�zի2���������|%��;U3�������������ۜ�Q���m��sd�QۥLN��[���ҫp�,z9���l��MR�h������1�K�,~.GVjRb�l����� �̄'óAF�j$:T�;<�6X�s���W����W,Y*�G
cl�L춊����g�O̩
*���B.Ԑ�_�,2C#G������<�Ą@� c9�X��ʢ� LP�e��b�D���c���]6���>��Ol�
{O�e�����ԑ�鬀��/ǲ�9r������=���;rė���<ؙ��zg��nY��A��p�a�T�:�5~�9��b���.�E;�����W�-j�Q��3��('0/������� ����dFy��(q��w�v������o���F���Q����Q䚥�Q�5�K��W6o�|��S���!a 0�3�8#��I��[tCuU�����	�2h'D���p���ja\SƸ�b���9�=a�L���fi��놌�  �����0B��VO�s:$�#�L��(��ZL�!Gp�TF��L��q����7�1�9��������	�V��9ka�D��AH��`xb.���Aח�r6C�Q.��N�ˉ��ROFQl�Y�zV���v��6�F`�w$5'���<��z��ȤeД��2�G��2 ��W��%H���C���ny� &ܚ>*�SN���m���߶|_J��S���f�y�]u{����-:�����Ё1:.���ݗJ4��A� �@t��&�@e!@LGD{�����g�� a;���� ��_��E����#��֕n/�&���d�H	</� +tL)�����6˶�4�7�	�3�r���|�#�,_9F@�ikt�8�[���A�?���@�!��O��Osx���0&l=�~�!� ���w�3�atݵ�"ip��	�c�a< �w���k�ʹi��	��|>%�v!��y�(g|^�A�;v�P�n�t���Q��K���)���5�[~��uw�q����zXkֺ�����[��jz`)8����{;D�7�4���"�(�p7vh(�ݩ�;uA�c������9��>��W�V�	W4N h�����8"G�(���^���năB'�0l�PX�F�1�Q�_����!3e���o�g��2�
�<Ϫ���������8_�w�I��z-��;� ~��^7�o�+�№�ɵ,'�����p���?�=�FZ���N&qO��>\��MozӼ�<�~����0��'�����alOm�:����7d eҒ��|��w�ˋr	�9O���-]�G9�6R�,��^�[�@x�h��)�w&��pq0u��aus ���#��q��N?���s��<���5�0���� c�} ���+��vw�u��.�r�}[�w��9ǿ)|�����mGJ�ꕢ;�q�c-�Xi�� �����=��j[��O�
>$�����'Ot�aA�^zi>%^/>���x'a��a�D�7M�h�S_�E���l�)��wd�B�:���Y��:���y�[ޒc�9��,�S��L�B�����s$e������M���>��g�3E�0���z�	##`oN�E��{���afۺ�і� � l���7�Xwڅ �'��ڶ�@�����r�K6l��p�{��VP3���/@ ���Z� 
������eR^�cʽk�����0ꅻ��2acL
E��,�����)<��Q"S64M0��ו���F�TQ��������i�2>�z��B��MXu�yv4o@�mܓ�Q�P�����������/Lqnd�z%��Y���M������e�.��V�ݍ��H����as���� ?���̓�� C癉� zV����� �/|���$��~�_�'e��X�\��e�FNP��x�esPs.���Z{� �ddL�2X�p�R���.��g�qƶQ�b~pZ���7�{��;o�d�џ	G~�]u7��~S��v�0 �<ủu�
���S���;��;~�Cc 0����ig�`�w�V.g�3��Cc��I��θ�u	5Z�(�sm�=d�~��p�m�96���&<��3&���=�L�byY��=#X<qp����g?;����E&\�rw]ڊI?�vA\p�-b��vRʲ�@�2�6���^a�0er���9F�	����G>2ow��R^�-�ﬣX>b�#s�1�q��5»�6M��Q(�EmZ��kDy",�	�t� &���/��U����2[���Z��=����v76���Zٓ%`������J�c�k�ޣȾ�u�N9B}K@�5��0&�M&�p��H�x�f@6�������91��5�(7X�β���Ŏ;��
 Qޠ��� *���Y��9X������ d���� ��>�R��(j�N��J �����tz·5��Q���D��v2l�&����4��=�}r<���BR�;��@
�E[�ي \�+m�6d�!��'a���g2Yf�*F%$�E�*���]>A�ϯ��W�r�)�c3:�y�5�&o���AL��Z��
�$� ܝ�|�+�<R�I�n���N�Eᢻ!$���H:s���81' cp.���u�00\%��_��_�bp�Ӊ0NB{X�E�b[dg�9�Y�As�E����ɒ�D����Ʊ#PF�Mt������B������H g�yf�>�Iy�s�o� A>@X W"Xhb.��I�a�`;�vއ�b�+�㱄�!GD-1u��X�GT���g�-���@m�m�M� �d��0�'�m%4A��9ʤm���o��v�hH�� ��D�8����H���t��������HbJ������]�� |��/Y�c��與��0�l�{��[W.�N���I\;�n�t�ob�{nT�=N���ӊѐ�y_�E?�\Ɋs��jT�\�E1��b���#�.X�����ר{~��pbN�j��a�]��D�b���=��
��6�hA8ztN&�.����y���vz�Z�' #�������b]3P,�JF�MqON@��cT��n��X�e `b��퇁���֊ \�,�w�S����@��)}d697`���zaĸ����q1n��1@�xk0�f�&e�]B]����!%�9Qk���H�r���͛7_tꩧ�X��f a�3k�����ﾜ���D����{g_�Cݳ�a��h���}:�����j��0&�TV'��*q�Y+�K��K�cdE=�:���lK0�1.������jpAR�s��Nx�%�<(b�덢SzO���
/�0,�C��xQ�Pg��4`���d)��k��_	��Y��z�����;@�v
+���+%Y*�Y14[!��� ��N��z(��я~t�	��j���I�0:�y�hJJq��0�@38Q��-���9�F;pMV$���DB[uP���,�%�L��Gς�2QI&�G�&������}ǅ+�{�2������y��4��[*wR�\�����I�V'�:�<�Vnw�q�$/�
��o&�*�@�\�{��{3{zI�&�D��d�2���'�.ty&���ҁY�u�)�dŽeb1!T���E�w�f�����	1x�i�e�:7�M��1�î��w�Ȳ�w��璙��YR�ַ�53,~0p��0a��v�#�EpU�pr���dH䃞�`�nɵ-�sB����wK��e�,�!Ә��� �P����l��	�"���a�{���/�\�R`�N@�� �0���^i��IV�Q�ʈ��<�fFك�x,��wu�hoJ�@XFo"F3��\2�'�]�s%�+����磤R��H�zR |��͛/>� ,3E�貔V�}�4��\�䀵
����I�v)e�&�H�q����ie���S���Z����P��*ai�(�`? D�Ȅ� l�f9)#?��w�x#t���5��X���k6(uS!g��$�J���X���~@c2t�g@��{B�`5�ıL�8b�j�Q��<h��6m���O���~��3�p�,���gC�ޑ{��@�7,�{�"Pdi�8�� ��g���F����8�F#����q�!�D�VV�#��aA��A�:�^��#|�E��BC�U6
%�%�� j=b�Lގ�fc��v�-��ǹ�؆��͹A7����=~	G��:� |���ޣ҄�j�0�vW�7�r%�sY95a�N�u��*��\��.�J�J	�픺l���J�fbq��u=v���iPf�k�u��s�9#t}�������P�<��2��������s�=FP�ɢ�s d�5���\���ʬ�	�� �`����������5�&y�8�Ir<	'�;N��=����H;7:��td<��;qT��Ǆ����e��´1e�A�|G2(��y�����[z�ߜ'���Ǆa�k�x�`D�(��ނ^	�h�
!��KY��r�D�$G�������A4z�=Iw��2^c�9`�|ꌗsD�� ��R�t�[��֋O;���E�}A����[9�m˥��c ��Ċf .������ۨTS�\jͤ��z���U�ͥ���j��R�6ݪ��ک�.��c�fsY��^S�7V�z}��j-�t�Sc)��J�TM�TB�贲�� > &L�ct���/كF?�yR�mW1a ��LP��bd�fň`j$����0��)���f�ê�P�� �b�ѠF?� <��t�g�m�E���a����ׅ��ѝ�Y�����,��5�r{?����[zP���_?�L���y'�9�Aa���rϵy������d�9�LX��!���_�F?��p�~؛Ǒ!�&���'�<ϼ�&H��p�$h3�.H9鷐&���N�T�ߍz�9��c�)��ฟvUl�C��o�d��;фd�M�z3W�X*�����J�Ԭ�{R�wn|�����MscS7�'&��T���6Y�ٮ�ʹS�\i�&J�63	�+�����ޣ�ssO*��=��nWm��U���j��J\�ԕ'F�$��\Q���?��Og��I�/��8AӑV���NZE:SV���w��Y �(p��>�:�VC�]B�Ыђ18����Q:���֋L�2z�/���(.�1M�ɐ"���m�l{�e�꿾`�C�*G ���w�Ű��ʄ�7��A��0<@�d&LPCꢎ����Ya�c�鉆pBU ���٣��,�~ �@v@�brv�&̱ڇz���ԍ���^��� ��7e�c`�����AYf=���r�|ݦM�^��L��0��#R/��*����oj��Vj����3c�2�l�w[+W�C{j��Y>v��욙�������l���}�n��YY�L?��灧����(��i���q����J�N3�6�r��A�A �+�8�!Q���vt��F�㊑ZQ�R��+NRq:h42��������t��R>@�c�"tQ��%�<;�2�RM���#��Rl]�y츑!Z����o����έ{�K�ee~�{�s�m��@AX��>�iX��,�\x> ��:wlìuF�D&��h�L&DT�$S/z%�����`)��S3p��})�3� 9"�Dz�1W2�0�)e��[.p�D�µ�b��X�QZ�m|؁pK+u2�e�-�j�����Z}nrrkk���[��k�+�];��� C���sL{����v�|Nm��?9>��G&���ƚ�R�MN��#h�0#�E������w &��$KQ��;V�
V���t�4ѫe5�R��</�	a'k�+�RcVC�%)�𷱿$>gԃcdIԝ�9v��,���<����@A�瓝Y/� �?�`��	�3�fT���E&,k\���sBNonX�h�1�@�a����)<��A �|��^{2���h6���Ɣj"Qq��;X9��0�&��M&�aÆ�O?��{c/5��a]W�8Ƌ>8�e3��TN��DjW&��Junz�����U_k�\���cn��导c1�*{��k�֤��k;����};�;���g-k6�[֛�sqGδ������R'�zr�Y�Z��7y�n�����1���*�#'��D���iH-����$,� �� �l�D�;����Aȴq�H���Ag�I6�:`��"���@eaN�EmW�Q[t'רC:��2�������v�(�Y���eT{>P��� L����'?9�6��N�pϨa� ��aϩg!;�͌���0�{�8^ ؊9����Fn�G����w�oQ��;�x�T����<��?�	�Q[R~�;�xE���eMxes����!�{��H�r+5R3U:ci��2ͦ�{VL�6�f�[��]��1kn��4�5䨿�D�����{w\���Ϙ��[1^n�N��J�VjW:�A^��,���8��	'��9�4^��R����j"|�۷��]�y>�0��D��J���غ�46Q0�h���,�`���t,�����Дy�A��=�fmٸ�Z,���ۿ=����]��g"K^�u�c��.�o�狃���<��|�8���\�B�a'ƬdQ�����`W䦀չ��kz��e<�4 L�.��zأm�u�V�G\5�g=��*:��qo~繹 <L�o8X���L�)C���}j1vd��k&t�&��67�sD��y��{D���.���Oz7�����p���So�;kd�4�\��j��i��>�N�vܳ~�����zm�?��/ݷ�وv�c/{׉+v=�S�������?eyj./��R�B��f.�xg"��Ĺ��t��Ǥ��>+���X.�fi,����H��ܔ+C�m�p ��  �Ah&=hPFm&���=o GM���T��I8��2�  ��"WL��F6�� t�I����l���΋�శ}8~�7x�g�,����3~����j.֐-F���ڪ� `eY7;�,� 4�5�19�Xr�m�\k!���>��e��c��q/z<�����(�T@�6����C���84D��I�e�<���LDr�����3�YP��>t��҄#I`��J�r�[���2nV�	�ҷKS��9�5=��o�?z��\��l�����4��������{�}I��/XU�?�֜��߲�I��zf�0��]&�0��t�G>�'$��Ս�8S<�9�L_7FL�.�/��Ĝ�ј�)���?��?�,���.ai�u��0�0����1�W����y�%�X�Łf1 ���C���!Vv�le>G����$.3e�! ,� 
�w�w�k��q�@X ��q�#�u���X^m,�v;�G�_�d� h��I{��/}i�&��	pрIlO�RJ�@�X&'m��<��B��2�,޹���t:��箾���<�IOZ�dµ[���vl}���C�0 �3�U�i�9���c���=�c;O\����E����Sˡ    IDATuO���g�����w���ܞ�k�Vfó��J-䈉�x�� �1I���K�v�ַ��uV;L�C��#s�7�1\:�
�$�"�������&��w�+殺�̘.���1�����}�p�ا��� v"ʮ����-/E���^*-ulb�&7Dͽ8��"G�Ar,2.�9)�"��f��d &�ꫯ��a�N8�	�_��_���ш����)��@��E�������ZFuv�.e/ًԦH��	�n�5��3�]2�'M��wd�`�Oo��Qn=������yQ��7(?��uѫ�F�\���͛_��'?y�bl�@\�L�����̊�U?�����w\���`�}Ҧ.�=p�oMn�����=O��'+�v֨����X*�K���Ǆ3�k¬�۽����.ơE�"�L��;'2��8�AV����a59�.$@�}��&���4��t�a,8@�$�u��`i� 1LV�N�*;n�$�����8�?G�T�81����O|"���Q��y��8]H@N&� s�pm[$��l��F�j!9�p#R<&b�4��T\%���s6��jχ'lzMm�� �a˖�3\���Nˀ�4!�'�F���d��U������?�R���96�E�V�}vÆ�}�S�z�blv�&|�^�~���1�Fy.'`o��Sg�q[��{�Gw�]s���z�m�)����+�����tѲ���c͙��R'5K�y&�E��?=99rX01���5BfE	�2{�����(�N�ڀ8��!�Æ��"󛱔�� 7 Lg�%"���Bg��$t@����7��ܗe� :PM�_��A�p�a�׏�.F������u5�{���|�DD `$��%�6_a+L�E��k-���Uc�vŤ��7֕2	�c[\C@D��w�7`��`�b��=J@�rp<�g>����lX��; �@F��,V�Nd�>�&#k
v�R���ƍ_w0@����c�s�p�6-k�֝��{�9q��z���nԇ_����ZsԶ��M�}׹��{l<�K�k����m��]��DG�Kt�**y�vޝ��|��&�F,S�9Y���@c������ʯ�J�<�){n?�:2\-:.�K�q��=0a�4sNx�X��v���\��\�t'6��	�vu9�b��R��b���������mʅ��>`	p�l�� `NbE��u�Ġa�F^l<&l���@*d5Rx��a#8�	'�'�&�]�;֏�� ��&�0���MS%�]=�kRâ#�?�  a����Rٖ��x>=Fۓ��n)R�0O�� ���/��u��~����Q��<uPm�+��Єg˕�_w����?;}�	��c�E���n1�{�M�NW�?�����w��̩V}Y�4����I���p��/��3���cn�@;;�Fvg09����d"֗s\ygG� l���ς�7,�侔A���PF:2�� V��z���5!G o8��/�����l����\������&lG��]����8]��O����*1ۈv��`��9`'��� ���Rmu���(��?+:�Sb$�ep���\ĳ�l�76�A�9S 4���3�F��`�7eP�Xj�� LY�YڌVN{��K6��L� ��\�n���l�0 ����]�nH����������2&x�
~�����۷^\�v�]�G�*�6S��]B]��4ӣN~T:��3�X���������ǚ�UG$؁U`$]ѭd('��e�'ٶ�`�%F���L��c�9	;����G�e�^G��xc7���J�e�Pf��06�}(�0H��8���a5�خ�\�Q�})�sr�:������N��8qE�Xǃ���; �$��cӡ�Wd
0�:� ��[̑A,9�n�),�KԌ��
���@Oe�����2p��;@��q��s�OAI��I�H�-A]����b�Z�qP�+��"gt��w��kq t,u��9�6p^E�W�s�R�37n|��1�Em���,�0�]�Zz`�q�O���n���_��Qz��9eӻ3q����ݵ�7�7gO�V�v��*�+�Jn�N:!��ſ��kci|l,5���j]]�����t؅Ҁ�vtB�	��N��g=+O�D�Mfg��}��N':�M]�T����ݡ�/���� 	�����$���;`QtD���#�-Ĳ�E���ܶ�2�DPv T�z?�C���	{ �� Y�20��F���E�=�A���u�Yy~ ;�z���xGdA�{l���2O��J̮I�)�ڪ��种aĬ�ע���I�r��B���Dw�(��+��Ю%/��mذ!/��_�lk��#y5�����O�9�x~�՚+�˟ްa�	�2L���X{��G�~n����o�C/�1������;Ϛ����V4�>�Rn�Z�.�M*�N'<��.��rs�T���z��#� ]���^0�=s�J��b3�Z��h)c��#G��e�E0.���_��.�!��+�`5,��ED��H�9l���ʈu�`HLb�"u��bp�]�]��n���^d\��@�+S�z!����ds�>�%�� f�2<!@�A�$P֫�>mړ6 �hK ���Cޠ]yw�Rcܱ=mM�<���x��F}p.�b����N,bC������g	��\��B
EG80�\�_~�<�>T2���y�	K�[�"��������=�3��=v�-��z�Rt��^�ɿ���[~k��[^����G�*�Z�=�J���d��M��	?rb:󬗤j��*$���f��r���KC���e��x���
`�A0J�2�	�+�As�	{� ���ɒ��눎�B�saU�J�ɽ`($����` �a��2E�Ƚ�Xb�/A��8�q�g�}��f�e8�m�Cu|�m H�h�<�̗�$܊�>�'[Vo'��m@���H7���w���Æ�x9�c[��@�bsM��͔���[@S2��|HD�@d��v�_<��7�$F9����IN��v��="�a�0w���;8�=�u.x+ō'��6dY%6�;�$�	\�1?�i��A�l�����+����@��91��y�c>=��Qn~��YhZ��'m�n����dٖ[/[37}R�2Smw�R���*>�7�H'������Zᩉ��nv'��v{>�A����LBi �u�d�z����,�
�-��he��	�z)�b�iuDϧ̰6�Z����T��6��(L�g��`��ι��cȖ�*?;�3�I��I��2���D�������$D� ~�^�=Wtw�`�\�kB,���"�]��U� );k ¬zd�מ�� °W��6x&�Źh�xI��sh�N'��=�kڦ*�I6԰9VJπ��EM�kEF���xuf�}��x�����xhw�8�����ڰa��L����}B��{����ǟt��xMw�C�z�5�Ԧo�q֪-��Κ�=?2V�)Ä�U�J*��S���ؓ�����Y�@�hu��;�C`��>2R*�	;Y�F+@�M\�'� G���9�s�F�� ���r��������\�9@�8Sadh��f�j{ ;��E|%�q}&��0�v�������E�+ھ��n`<�yœ�~aꌥ耰��;yw�F�$t��/�b �=�7���t�#���jK@��L�~͹N��,�/�2^刮u���|~���}D	�ߌv��&.�G�C�6�]{��0����b���mګ�Vh��W��a�]��kN�������M������~����7^ݲ����l�t���*ө1¥4Y���N>!�uΙ�����R��������D�B�U��#��QtⅲEw����7���_W>>׏�8~.��,�w9�spY��5�% LP?���� "�ᚬ,lqy�g&FW�]3"��@,��Eh�H*`����3��������, ��F$�����6n�-Ѿ�%>Äq�ѓiC�Y��xC�O.�0LM�g6O�A����,���n=em���>���q��'��O��T�2�~:L�L�v*��se����(Ca��1�uw�y����1�R3�aQkV�s����kl��c����~�c7������<���󸍟Z9���WOn���k�{���S�5��6Wf��&'��U�צg��ϤR��N:�Ĵlr*���lwC��H\��]��6�52B�#)�����t�x|�C�]+v��Y��;:'1���V�	���9�������6��� 9�DB����;�%>�%�ΚG�x8�0ug�u��8�s���۫V��N�2t�Q�G �� L�	_�"�ri�G�6�d�6�@�k��6��b�y��QF3�2������a���Mm�gs���c]x��z��uE�NC������hO��>�ܴS`��!����3����}n~��z	����ʭ7\�~��W�g�n���I����\J�j����c�g��������L%v};���n|��m[ߘ��e�S�z*7fR���J�R����������/����Dj�Y���E�*�a��
��#D�#��{a�t
2_ѱ�p�C/�r�O�C+Pv▉��;�0 Ё	Q�3"W�v��vG}��g�	����/oT�ڟ�^�sd[2E�ⲛ �v�	�c�|T�Q2�����I `r��	S ��O7��m3@��e���@ȵ����=��1��,,bGp�+��8pM�E��j�� '�%(�;.tr��fH@,>��y�������D!�C�0�h�K����
��6�'3E�"`�\�Z���_�t!jh�v\��	��@��Z�j�S�J�LuC��?:}Բ����,j��RT�3����*w�������dgv�T�����Tnv�7�6t���T�=�ݗ&''�o�Ư�����nTD���F�F��AX�(~�;'P����P���x̀����
H=D���Pnf�)�g���Â���0/_��R�C&���D��sd& <�	kqp;��;��j���y3���] 󐛁�u��~ G/	ǐw���c�##�g,�׊R��b�ݐ[�I��3���(_p'yv�KYB�r�w�Q;v~������}�h�E�1��z���Qtnq�2��ā��Bl���~Ll�T�@c�Z�N��Ax�ƍo\��7^�v��� <3τ��~�<��Ԗ��<��/׏>������~ ��s�����o��_��{ǅ�=;�9Ѯ�f=3aB�J�Z��ȧ\M��qg�Uӹ瞝�y�O�Nj�z�;����1�+���;��E ׵uFZ�HqcqAa����袟;� �Ɓ�c�0��U�ݠ'�iGaY���+��޸V8���; ���s�L��zǮ���A��G$t!2aT�`��?�Êڃ	S�)F�X�~�b�c9�,�XO��9�- ��}�ss��f��}��)�xM����jM��R� ��sb��A��#�0@�����e���}����"��������9�������3E���6����M�ް� <vˍ��ٶ��T�M�R+U��t�R%͕ʩ^kͭ\�O�cOx���1_��Mu����~��'/�}�'w�󋝙ݏK�4�棭z��]�N%�����t˖�R�\J/;���'��͹41�l> �  ��y��0�;@d�<"F�v�^d]	�h���^l'�W�2�8����K�,aP>�r�atb\�Q�4T���L���Cd�����!0���EX.@';Q��B˄s��b_���= as���xG ƞG�Y�����߂�e3l,��`ɮ/l �m�`	pAg��F�oT�+%6Wͩ�82Yȹ6�AqQ�����0��*):!�)N�.��/��{�֕OH4�8@��AC? ��c��{�ڻ�]�����N���V7�D�r'uj���Z��}ԉ�j�#�����q)*e�56m*�X{�s��|�-�����R�������ިݚaX0Ӫc���'�����87����f�����w�`x��4��|\DA��ȋ���p#iB�<���X`Gh Lg�?/u��ϻ��������bd�0�1�c��t5����3 �V8F�c�Ja�_�n��P��.�l@���o��
�r8����w�3��Q^�+�6��K|,@(�.L>��m�u5_�-F���W�qxs�.G(��<�9y��*�%�u�,�n/��A�Xy��+&�)3 N���R�0\l3 c�\����p@Y���i�Ub%�_�u��z��z?�L�+�n����۶]��5}T�<�zk�E���DoM�ԩ�ӞT�4W���1'�oj��?��i�൜�X�cN����s�+�����s{�����i�*��ޖ�r�������4��ؖ���ү��/�S~�������T��r�8p=�d#b"K�E�sa$�0l#f����0��lh��ha4*߹-����u�`	�8@P$J]�w���N�ŉ�~Unǖ���Z'/�R�	��9�C��d��T^B0���vڼy���/ �<Y�-��}�M�CzDX1vc��h�zbf5�q��=����a�������zl[%.]Xo��)#�xõ���ye����9 ��C<��;����q�xe�{��>Pd���6�&�LD䏃L|�Ŵ��F/�߽�D�����eC@��0�,�T� �ϲ;o�t����hͮ�g2��[ޭ���RJ�R'ͥj�WW�gc�1�8��{Ձmq?�2����o�8�z�֋V��E+ZӵJ��ʬSn��'���c���.u���8:�Fz�ǥ��n��f����Ra!�(3���� \ԋl@����߲#����1)��VL�=��8 j�"���� � �	#IP&�W4�Q@�q�Ƽ����c*up>L���fۑ������(�Q-h�HGqr�g��mڴ)�2���d¸� :� ��&�8��.S.z'�_��O�m�Uk~�{�.n��GD Ҵ#�y�l��[d�܇Հ���p��v��l`㑈p=nX���_"�������m�6('�}'!x,���(C�] s*�͛7�aɶ7z���;jj��oZ����Z՘>�S�)Gnj�rj |��4��33�������cW���\p�(F��c�������<�����wl��W5�{��TO9�|��:�	�%n/U���N'M��R�>�M��jtݤ6�]@Ɛ^��e����Fo'���0V/��wq�.v נ/��	�zq��� �!U�%h�<#:�0&A�c�dγ��I
�B��Aw�ו>��;���#�At.�lLP���>�腗���W�` ������h��!u�{n� ����Ł3���A5�Y�0n��,�d�X~���|t%\tã�CS�y��(\5ʻ�2�z0�D&\x�eH 1"����A62*Sv���>�<�F��\�h=t~��>pRe�7��s��Ww�M��Z�]�r�L��f��j*�}|���Tk;��]�͹G�'�=��;^��~^w]�7l��t�g�߽������_&K�&�i�!�d�x�>�l��Ff�,��Ɲ�q��1�9�>�H�+��ҹ�4�� �я�c�, �L�bXLܙ~���\����OC;�w�S�I�{�b�5v�CY���Z�r �&��:z4����;c�A�:�SP� laYx&HD֓��^H�_�3:VoF�6����w�!^#�Ɂ*��L�+tRz��XV �]H��9Q��F��
�Q��Y�{�6{�a���8���$[��/���x�ٜ��� N��%�����_���-7�κ�;^��5s<q©=;�0aA�=�J�r�-�Ӯ��={V��������>��k[�,����������2q����w�󧦧?ٜ��`���"W(;� ��w��<Jw�	�J7�%��l1�Wt��_�A0C��E�l)�1׈/��|3^��b����͡;6;	D�0 �s�j.�'���)2�����s2��[1Z�/����f��p2v�A���k�J�  �IDATtQ�!u����"��4�5f{��V�c�@l�5��kjkʆ 0�a둡GV�5�������`��s,:=K��đW /�d��=)c������%K����ౝ��^���m/\՜9�]�M�v=U�K��.WR�Y��N���s�D��k�jc����������f�66$�tC��M�R@v�"�&2J?ը��q*hq��GU�6?Z	!T�(M?�&�*�
��T�U�4���!�/0^���̽��9羳g��ݵw�����̽�|��9�y��u�4SH�^���]s���6�۾Y��\ɩ���_o럟8�.^xP�_��?����u��8���BKA �q�тf,;+��t�@|Ǫc$a�lȓDH�C1P� �������Z�� L�<���!#)��]k�׆.=�	�9b�G�y��#w ������Z�C��]�����[�TSDK��-��3��N	���#�7���I��[�:�A�.��~��F>(����o+�F~DŭF_�lJ ��?�j�C���<=|5�Cz�vp���P�����B	=8�SY��5�[3I��v���g���?�	�<cn��+[��=����:ώ6ϸ��P3Ƚ��6�`:����,��@��\ԛ�zN��ު���,����G�vKc�TV����f�>M\z�M|tW�^�� �c��u����C&)؂k
�v&o	[��XNF`R@��gu@�5�_��MGd���I�A���݈ &�x�� �6M� ���@���D-4R6�H4C�Ǯ~�^��	�A�a4B��$)�r4�$��E��o�k*�@G�^}�U����y�\k �A�W� �)@���I/�2�w�JI��m��,=P� o�7�s�<2r#�����>�.�G|	���0ʄ'���pA;F:=�oS��	!&�'���?ڷo��o�Z��Ov杧�?����3�^e�Yd����M�1%{�g�����3�gU�����~�7��w�wYe�_�rx6)�LM�p��or����1�llL�f���]��ӫ��z��LN�U����hvz4Lj�%�0$,��L'��T�I��'�� `��I���#�`R3I�؊��.�`�F�du�����#�L2�0|a����(Y��?���э�ɠh��&�FPG���b��cF9�� -� �>�`���/�0��� ��$y�-�݂W���n�s��'�A;��yi�`�A:a���6����3�`��Z�.�v�$�?��0<S���;T���qz9vA�3 c3�%�K�w-���������_�+��:K�0��d�G�qݹs��W����\$y�z`��;	$O�m�Hpɐ�A&��ix��sΦ�d�R)�a��
�t}���I9<���=�K1d����?���ĮQ��j�M�PZ�F�R�ګ5ZĪjU��Ԫ��R�����V5�ؔ�����γ�z�s�3]��p��i��L�0�zo�y)@TYfvf��LS"-zDm�0z�EJ�Ę�y0P^�3�����=s�C["	��sPD8#���ﾶ�|B�����o��'	w��
�	.�S�<r�qҟ!��&�Rf?i��	��\�Y�N�mO�	$v��ģ�bHj���qE�ʉX�T�($E~���8�kq��~��s��~��VǈQY0�<��wm�3n�*e(��!2Xp)W(^FYȏ�M���ڐ0z��(���1%��Zp�À&�N�[���U�rZ��1�Y-E����X�:�%����Aio��ޘc&��g�����w?Ek��8�-�6[����j�1����?6ٞjW+E��M��q�F�I�6���F2�����D�< ��D?��������+)��n8E�	*�������V�m*����2/��}���$Q�� �+!���6h�I�5?E,�qI�Ʊ�6�:e���� Ì䠀u.n(=�f.oZ�*��ڌ��tZ�O��.x�*uS�ʩdKҔx+��$��ðc����:�ԸK�,��M� \����5(��k����wh�l��h�m��"�Κ-�Sڱ/�G�,{}!����;�~���T]��q��\���o�X!rB�:A~AǮ�w�ґ~k�D�"%ᭉl�4Ց[�<����3�XGP���:��[<��|^�8;�0�&g�7�K��8��B�w�n���aEߝey>�o4��v��%��4D�e�~Ʊ��?Ӿ�CM�5y��w�k�3�����d��%�G�o�=d�;���I��<�G N���v��<������0n�S����'� j���"�C~�Ñϓ(�<�+m�z���{@I���pY��9�qʇ
�#��O|n!�}�T"[��*yy�Z3�g�f�
����<��>�!Y�CF�����&Gk�sX�yy-®����2vW?-�ʁ����g���,x/F0��H��"Ax�Qu�����?�R-��p[�<���1�\�Քۡn�G�f�d�%���{�𞙅aF i��qee��#7� ��3��׏7���;$��iX�z}:��`�����LuB��?���<��("���y_���[9��ED��\�P��Q_!H���I���B-���M�B3jf�={�F,�7j�I�6	)�8�_V����>[����wkZiͨ+D3#�0��0���o��?��y�Ʃ7����?�?�:�>_��~�����Wn�J$����-�y�w-�U�!7�=�K���62���U�f��7	���	��I|���*,-�\eF�I�G��Q��x�銃� ���}�tW�B�� я�<�.s�վԣZ0y;�pE1��±G]�x~�s��duF1�T7�N\P�����K*�d�5H5��{���៏�d'O>���͎���xr�&�{�կ�B�;]Iwȷ�*{���Nŭ? Ѧ�Y�6���5Ɩ���Z�g�n�M���d��������̈́�+���]�&Fܣ3��ȝ����\��m�����J%�7�N.V^���lOI�W`��Ԛ�;��rFM�hO��&kSkwK�F�d*�=���e�yU�2J�~��s�<�<�m$�ȁb��A����F�1$�JCzG�9�0�X��=@��L\j��nl�˓�7��d��4�̈́���=E@���Y�����Y_ވ�o��N?�vҖ#b	�
�{�� %�R�o�l��u�i3����7�( �0_#G����W:�z�F�I�Sh�_���Ĵ-k	y�E����uh|�wrn�I���K]���+ԥU)�~��J�M��h:��,���0XyO0a��W�m����m�	i[p��������b�w,wk�n�i���2���|Q�aӿcOd�����ޟܟaP[_�BV!�,��
���I��ʠ�5W� �>���O1*��T��C�".C��±�$��&�^�o,k���`>������b�=`"���r�ʼ�"���T����n��րj�����B�������!�������Ѧ���C����I�ǯ���>ZHc�K�V��
�;	�`"���X
���/�����$�Ďv,�[��5�8��f!�-F�[i^�G��b�#�ۣBb?B�/_ɋݭК�Gb��xI�ݩ+��@0Z0c��]X�)��"����lps�lU֩ʑV
�&,��焾��;�E��sx�g�k���=���qH��/z	B�=���@�!7l���������Y��K��WCNC]�����:�0�w��0����ɻ	�%�e�4��()��c��+iY��l!{8� �j���%�&�Z0��ә�<���Pf��36?�[�z0�M�?���x~[�੓I[*�" ���.�$z��Y��f!1����>�g���D��UgΔ��2%z_�ֹ�\
���82�~Mg�kTZo�%s1�ˑ������ݣNw-��)k1��o�Z�F&WК����D���i�5j��W���r�mEwm;�u�`��IP����P㕗~��Ka����B0�A�q&�>B.���0בTI4K�� �i�?�R��1u�03<ԏX�7�˂%'�mj�9h���^����ivJ��A�P�4R�m^���P�MݸY��� 	3�ܩ��^	���E1�5� ��$q��lJ�O_&64��%*�����b���G��O�w��;�����F8P��cfpBiN�-1R<0#-p"ϲ���R��,���a�F��IO�sd���e3����I�F�]&�N��74}$x{L��*۸9��ԃsNVق>����{6�k�9�2���[չ��y�0�H�e�UKGd�V�)��
�?�R�:���l���<XIZ����l�j����A�h���r�W��y�8�X�;��쎈~�)S�v�O!��ێ}. �B���t&�Y��)zG�A�2y�Ÿ�3y�`�
��PeuW��.�id�sĻ���r������!?j�6�#ي�V��}�;�v��#7� �eqe=��q-MgDbc�,����<�=��]79r˫2���x3�ȧP=���}���u#AQ+��|��CQ}�Qűq�E���Ȳ� V.Y`�F4���w��o��{@���x>��	t�@h��;KmO+K�ҷR+��6,.��+2c��A����-r	��Y�����WZ,c�����2�*���1ۤJp�����h�J�������Z@�8�/ILM�����W�#�'�����J�|����q��ٱtǀ���Ϸ9��wW�wB�B�lk?%���������Κ�ꨭ5 �_R�F��Ԯ}�3�"��'?�2�S�t���(>����Ν�O��\��p2Z����4h~{{��8Z>��#@�Πu�Π�S0�.���sF	Pԭ��d��H��=��PX��x�v��o9q���="�J��[P����{ǭ����;o���NՄ�6��.��mE�������Ҩ(���<�պ�?	~�W�-e-6.�$���ɋFaZZ���?Ǜ������cU���!r��鐵�����ʗ;^';0i9fI���i=XI��ɝ���:��^�\�n�{7��>Ԋk�����>�;��Z_���0�7(penHV�3�Sx:�Ҹo�<��{@A�4�t,r�A���hqb�&�au=��S��
��.��E!��;\�(l
R�Tݖ�V�^�h����Qt{J�~aulM1��Z�'�}��:��~ϝz���I��`�ϊ<O�.��GS�؜��i���{�k��	�;�j���\�Դڹ�,`��>}M�=;?֘����D�bZ��"��V�aH=��ov��,w�pn�ө�o�Q�+�/?$U䴐�^��g�:ںf�c�j��д^�w'2�_�&.F�m8�z=E�T��|�����^�*`���r��.H|):�F0�ޟ��_�2���2B;���P�D�	��3�'y̭]]CGmIR�����B�|v^�=�}	�߯��5��M}�XI���n���2�S��ToO����ޖ��_E����KPɸ����Im���ˊp���D�l�"G�,cC_���G���)��ui|ۯ�u4�Q@N��)j��3�7zœu
���hPۋ������|�q-#&�1E�vK��/j�ET
#���A멃�,*-^�!��GA��T*u�*��+�6�6PŁ���\e4�Ҕd���x益�������m��Bj"�7.��̗m71�!��U����;<��o�]�K˰�u������������񏯣�S��FB��tC�_WW/鳇Z_� Ps��k�Ѝ��x �����ö�nv@9��s.ƒ�d�������%��V�C"��Y��n�qX�6�G�?��n���$>�z�c��,� �WF�.��}1�{����
W�+g�VK�Kb��6����w:Z�%�Ko\(�[�s���������2��=��($T���.q��hB�@3%��]d��a~~GIɿ$�Y����������k�*�[?Ceg�3��rƔ2��v���ގTڵ`�M�oOl��PK   8f�Xt`�,s ʉ /   images/94a69387-ae01-476e-9716-f0367b107947.png�eTTo�?:4��J	��4H��0��Hww���1!!�HJ����ݒR��1t	#R#}�������/�Z��➵\fγ�����s��ik*QQ0S�@ *�Ǻ 	"�#'>�%q�#�x��O\/ɟ���U6� �n|��#�p��>��`����n�n���B/�<lm�vB�����R� ;H屜�w��Y���F��g��w�?m׼H��TaU��I�^i�"��F��͸oz�q��q5n��\��I�{��hU�oU����.VL[�S�yꒊ��H��(��V�r���4�G̶�{b\�ӆN�έ'�;�5NŇ����^k����e����� Q��}~Uv��3���h���ʠ��\ʀ���e'�����3���6���'��2�����2�M�TM��HH��ykfK_t�v|ġ�����.�干�+�_��ɢ$�Ұ�����|2�jN�d;��[&����aMS���*{��|��J	�n�)}{�r{V�z��>�����k�uu�Y[NfB�\�\:������S~7�����Wh���3�\��()����5BR�n��G�3�l���l���u�%������������k�c���éb�޲d1��'#�!3����룓�Oɕ�g�<��7�mB��
z�]��N�`�;13�S�
�XE����.�L���x�DK�=6��p��[||s���+b���Z�W�q��wo���>��˂��ӝS��l�mW��黦w�}C�J݁p��x݃�����*o~\)�;��m���4�׫g�+p�?с����<��
��n�A(7��^��*��|�U�TkT���p�&������9}�~Ʋ��@�E.,�Ta�R�i%p��DS�8B�=�21|<3��d6��;@U�{ �H��F��(̫�r��K�_����w���QT�q慧����O��t�f�U�i$����KKO~�|�e�O޲3�U�칗���������Mœ]OOך�x��`��t���2���1��:�}�ޜ?�����&�ˆ�ٷ.�4�'�+��6��&��j1��6FjY�k63ly���EƤ��\�[M���0d���v�TP��K,g��d�D%.�},�k����P�W_=��v*�pr��Z�]��Z뻱Ì�˹�W��
y s�\�&.n*x�ج7w���H�G�<l~;^�a;ϊ}�˜.��'�wL��jx;J�.��h��df��r ���jt��9�\+Y�@��9�oxlť�`|`�%/�?GC�M�[�� ��CWaXBUTk����Yڿc���j�\�@b�v��f��C��_7�������(�����Q�to��*��֪�:"x<鰽>_%�6�[2]M�.}�u�65i��0t{"���3��o��ף��!gzt(b�s�f64����|�G��P���93^e�$��R�E�|�F������4�	QCN����ab�+QWoQ��68�b�j]��[R�Ɩs��p�j�8��?�k9�����Cfdv3BN��g�S_T��2�X%���F{�"���J%�ib�{# qe��{����[�3y�������3�K���ٰ4m�>a\���#!zd�h�V�P��/.���rU��T�*��n��;Q%e��C ����A��щ�E
쬃Ƅ�@��}�qzNh��s�d�?X��ō�p5��[k\N�����O�{���
���j�C���"ޙ-�^�>����N��	r�o�v'tj�Z�'��m�����cQ��u�I����W��fd_�n4e��yϝ!�.�0��[�O��a74{��+������-�����bX���Ň��(�R��u�K(����
ǳ��.��������������M��f[�M��kץ�ʨk�kqٛk����h�EJ�b�8a���Vsn��I�q��k˺��� �M�Uw;��:��SP����]���ߊ/ζ~��)�Z���-^0Q��	�𙓄ϼm�"SK�W[]Tϡ���+݃����%	����f��#�.��~_*P>,⢕� ;5��u��}Z�9`6e������L�u���/��P-�j-���
XS���掌tjB�m/�~��G߮�6�`w����9P2���<�V�&��X�z+<˻2�ܤ�$��ZT�G˲L��V���^�[}��4b� H@A�
j	&J@g�_��H����܉Ft漧3���p��X�od �hS����0�L�;̀��5��3�.bk��s *����`,�9۳4��yxx-f��%?E�!e<7�4�ck+~��D���p`u�Z����E�i��Q̈́R�]%k�bO�W�s�Tz�0&���QI�GF���7��k�������{ƅ��g����?�z}6���2��U�������L��ͳ)1*�ɘ�y�O��Ÿ��"����e!��B�0/� �^�J_���/bײG�|��l�g1��"��y���?����G��=}��{Uy1� ���# p]����ԕ�>̀k���{W\�Gu�k�+%�kJ;�W\���B�vndf
µ>gh�mρ�a�{�(4�$j���'#j�V�a�bX�x��v_m�z`��0R^��ǲ�w��`]�in��m�`���'R�-�?�����bTk��j��TP���⹙�̠f��.v��ڴ�F�ͳ͚�U��jqƷq�y���Pn6�xf�p��R�l�~}f�CL�T��#�:�#a���!;}ǯ*���IDZu�
C|���输�A�ݎU7��Y�$�63�Y�Ki�#�Z8���֩�p��eB&wt�Ou�z���Ź<y��U�@c�
H����#y�ku�z\%���D��S�&��_��r�yy�?"P')�R:N�f����~�b��S�;Z�g�j&UJ�H�r�a[��Zf3[��;śN�o�<��:RQ�ʏ���>�� ��K�ʸ���P�2���L�c4�e<21��,3m<>A�'F��Z}�%B�����dt�jy?n�_�@�3�k��h�F�|�Q����.�ovT^�2a �Jx�hC�\D��p_�@�/��#}�^�=��ǊHs�����!9S���!T��MT��������lR��o:��?Bڝ���zGk�P��7R/^�o|+����c;�`ie.;q�xO_u02�M3p���=k���(�ni\'�t��p��Z[� ������'�K*�M�l����(�%i���}Cr���rS��>�˳��̌d�~>V<�SIe%����|����*hD�.T`����晷c���MmD	�����m���8S^��z�k5��M��ŷ>ͦ�� J��eg\�C��+����`�������y�?�y��RU�[|�T�_X-	_T������%���7�kXLڶa�xC��6�r=ܕ�)���p������b�8�J\pj�j�����r��� NX?@z�d������ǂ4{Τ̯m���� �l5Q�D��|�z/r&!j�5PܰP�4�Kh#RW�`��=�J�l�@�� �j����$+��;+�2�	F����b�����u5n����y&�,T6���b����F�\�
���]a�z�3��2�CS��L�[�f�q.&�g�|��(��CeS��Y����^L��R�l(�*����5���O+�/�P
�	���.����ONB>�4�ff��Ϛ!=�Ԙ)q�m���8�P`t�Ÿ(��<�<*�$Jmx�.��.�!������aq�CF��a�  ?M�k���OC��wcf�l�.�yDKkGB!����vx��6��XHI�;	t5���rr�2�Χ���AS��4Y���r��/��4T �-q�zsi��w�4R5P�F����;g�����@?�s.`��p�#�
�)P�+	��Π��vi�+d�	�����:�9SR���cJ*�ue]S
\O#�K�W�k^��Zb��ҳ2�]��G؆�}�K$R�~�2�����gٚ�jVU�E왤U�.v�M)�:��`+�U<X��싃C?�������.�� PN�}����:Q�֮�Ȱ���4~��f8�T���}K���;���=�\��a�y�c .s�p݇�A��o,�N��7˳[ p�݇�> �/�E�]ҋ[��f�����h�������U�$��췟aXNhf�Vxc��,�p2g���0wX�Y6s'^{?	?�X��&��*�&������O�B�[+n�{>��gG���|\�#l�
�)��*~G�Ʈ� �C��w��f� =��T�[Ş!lK	�[���4���뉔/*�99K!|��D"��ޜ�����M�I9p�7fu~�Fq��։٧�MN�AE-�&8%4�#�ӛx& �-a��&��;O�8}0�W����}h��I�t_��u\3Si�M"�>�� `V�:����Q�<)}��ӈ�PH
i���
�.k	������u	� �u��g�](�+������o���Y��1:��XNҘ�b<�`���T���=(��}����>�6�dv;�+����鞩.dD�z����)�(\h-L_-���)�-�Um�M %��BBu*'��m�	�{%�MCe]����9�F�Jz��4	�C�/�������+���� ��{1��j�5�hԁ�k?�|�ב�UJ�L�ky��V)��!2����雧���1�Rן���wz�����f��ɺ�Ȉx&6�-�P��M]
�@M{Z�m�)9t�Ȇ1d�2�6�LE�s�\3{�7�-�յ��?z��K�6����m�q����K���`ۥV9�������W'��4��q��Z���7@m��fA�\��{[�	����xZO4(�/�hh�	R�~Y/��$�D�ؐ3�֭0�6?�~	��Ĉ�s؞���V�3U+!��֏��Yw�|���F�>�V&�1�w�0��ZRj�d�}>��1��ւmj(���ʑ�ьCVF�2�������y� ��စ9�R��������^�u����赾�e��ƏSz�V�a�Y�7hu+Q���O��V�M-�0�t������-��Hpڱe�]mJ'T����*п�<��F�����6~���s=������bn߽���/{�-�8�:bԔ��S�C0}�C�Ԯ��o\��1O_Y�~]S�+a:>�s�T�2��z�Q���R;]G���ȿ����AHw8Cs2(p�	�y��
�&���D��
��<�z^��\9	 N(�(��2���-�>��	CEHv�oq�W�h�[�&�C
����VJGm���X)_�R��n�6��K&�~�Q,	�t�	�Ѧ�����Wv:b4�ד�h"��p����T,��I��ۛ�����H[v �oPOA� �����bT�ne�X_(�F��g��_x'QE��@e���;�#��G���4��T���� ��?L���x���fSN{,�t�Z���$����d9#:n�ZM:�	�v:o��_*�E��>�.=��GQ�^�@�V���`o��3��夿���z�ߑ8 ���(>��爬�Pm �R:%s� ��Go2vv�d���A����}�B:�����c3�Ja]���Q�:#��[�uy�J+�_{$�Q��;ƯU�~�qD,�48�ݖg��@ۃ	�c�/BaoM�)p}}@B u+�	���,UD��!���{25QЖ�ӑ[�B������7��{����Z|���Xm�@�`�ی:�q!(�Az��C�1�/M2EP�/��KMlj@@��G��8��(<6z�j����A�+�� 
���Jy�*�T�Cr���_T�M���N�'�lç��k4��hhnZ~K�HE"��u9���AA?�TnS
�3��.�4%���$#��7���ڋ2{
L^��U�ǄI!~ڷP� ڨf��<ܸ��!_���V���z�2?2=�l���VRL�d���ss�7+��	�bz����A�r����e�>O�Vh��}Ja�)W ;�����i�!@����N���qL-��a��L-^թ�i[D�a���ܧ̌���⊴�]v��A����lz�i?��e��B��؎K���MmD
�~V�!�� ��WN�ˆҨ �8�00e�d��w�(�X7��R�7ш�@9�>�-~�9"���'�{�h��a:1�@�qe���h"����uf�Y��p�c�`ɛ|��lq
\�M��o}�c���m^4�:ϻ/����C�Gz�W��W����j]��HRȑ/��.�'A�u��I�×Goʠ2d����|��m#n�rMZE��hڻ>��M�"��^�'����(9����i�Ēo0a�A�u���yt�����=W=�!���W��b�y�>~rr#h���6I"���ɻv���$N"̜ɌX{`��� W�SYH�	P8��I�Hɒ�2���\ӊo^�jo����ɝb(Y!��-vpj�t)��q�ѣ�na�EVU��������o��"A��}�*$��r�����rD�����#�� l�+,>�1a�/�����&(����g�+ñ�ܶ�ۜ�*�]�B�U+�+ 6�!�B({P���*BV��?1/ǹQǀH��2wJ�Cw��ca�{:��k����4����f���7dȿ��;��I:$xzZ�d��� ٣�<�r�ĩ' o�n��f�����G���
�쐅 x��PJ���äN��8Ji�[�K&'�����S{�re��� .F�V��L�%@@F�����t��"���c�<�+P )A��<z�EK�܂Kr�ږ��'�0� ��˗�E����>S�Il)8~ő�Î?W$�B���#�����=鰠GK�j����Y#Đ�9R�{~��K\tꤩ{���i�Of��AY9P! L���j	}, �O���= �:������Dp�Z��i�7Qʿ�Dc�$[�m�MH;�C0	"���F��o�I��X�}� ��|�
�<D���d_m.�5!�T�H�]��`�g��!�P�"$Qj�������հ7�:�9�Ҹ�l:�F�U܇�u W ��5� ��%ծ@�x6��[M4sa��g og
hD�,����1WG�J�1f��eS[--����Y8 �}�A�x&���[��9m�1
�<&E�2*v�u㩀眖����R�T�@�j$�aD��Х�Ό{�TMBz�
��-B��� 'ٽ�=D�.��^1ڸ'�o��h:E�Q�o��\�J�D���<� ���{�:ڑQ(��/���G�k��l,q�Ɂ&*�d�葯w���|}�*/�� fa���"HJ�P�
���3%��t��Rl|�^�8�7.���wf�:R{�w��`�9�p�F��H�����0A����3a�Oګ�M��Am[S���^���p7=�*I\�����.�ܿ�(@� �8#�yQ�}q�eDϛ�e�:������X�|�ϵ�b�.�ޡw:,<�s��	TAQ�ҷ#�	E�̸CRYh/Z���ġ��0��s�]�L%���H"kQڔ�8���R,2E�x�"~�ҿpg�:3hd�a���˹T��V&ֶXs:��P7�[b�+�!d
��3��x�3_�j�<���7⮞(��~s��?$�v�n���7��f������τ�OV�+�(T��@~�����Ѽ����}�;,����dYV�A˱��5�ܦM��`~���;C�珖����Qг�d� ��f�a�=:)�|�l�oz◓���pl�흽��#��d�RCv����^����_�y���KP�+��#�qx �c��eP�%Q�Z��ȗ����UT�.G�#"4*_b��jt�8a'9^l\���l\�a٩�==�lQSe��u��]ix��i����9Cۥy���Zזp��=�����(����;n�|�]�J���L�EL��.�by��/�
|�v�-���&Y����&Uջ6~d}ߜO�e<�|�&<wB�yW-
�0��/sF���7� Ͱ�^�=%�\:��������P`����^֥����U�!~��E쪕����31ƒ�6�ܮ³�o� ��S�^��Ui{I�����h�ГY�͊��>�����4��QZ��*��L���{��eJ����|4�|�J��<+�m.4�h��!�&b���S;tbr|�"�	�L��vj/�S�c6m������Ҹ�NH�sȞ�2Z k���B�ht��e5�����tb�~�/=����w�++��P�b4���y��(�E:�p{ñ��P�����iׅ�Ɛ�MAeh(q����^�c�� b�E,,��� ��|��
�Y�)<TI_yKT<N@�e�B&=m��끦 qv2,��|5}�d������
������LX����B � o�W!ZP/~A��jT��K�[�#l�i0���k`s
$t�Y�M�$�&j���i�oX�;\P�E��;d�d��y��/g�?H� �H�:Kç�5��vK�e>[QuvI���`5���"�C�5�r��m׽��Yo�*����$�γ��]S|��!JW��\H��c ���Q
�e��=�.�v����ATJ�J�-�O"�:7�{a ���`�V���2�K7�����:Q5�}'�xc�?��z�/��#-�F�ȍ��^���p-�~���q�I�} �aU�TM��B%�ǟ��՛!�O�_O&����f)��_��`�>���d�G�aRNoxV�jj����d������Ԩ��q1�jggH�x@�&8��m("�!��PNHl
B4�A�Qa;8�j�?h����p��2a�#�[�۠�瀏wU�JPLh���|��+�@	߰0kL�,�`�^R?��6^W֭i�d�Ǚ��B�~X��|2���j,6ӆ� �[�{�w�ݚ��I �V9�s������v���^�2C�a�����-����
���t���(�<�İ�H�m�3z��:?��l�Ҹ��@�N8�˶�_�+�x5���8�@\�A
k�&AF8 8��Y��^��+m�l���-ٚu��Ű�Ҿ\�"���[�!d�6q�4٪����T.���jKJ��U��:D弢M2���j^��J���@�4R�
3RV��Bl�|�g=����7D�M��� �
���,�S�
VgOҒ�PD=���1������V����|����O��,B�#W���|��������:�����AH��&�'�=� ������~Y�4�F��A�1d�|&��O��!ءî��k���:����Ȅ/G�K\���6s��5�#��]?��J�+I`�ۨ�s|t�%K��Ay;�B��
<Á���
G�};C��j �h�(�r�I���v�Ćw��v�C�֍�(P����A�u�z�.�ҟ�
c���!�$XA�Y��<���B��r��Ĝ�[?�P��Fjm�.|��rd����-�LOG�?�u��q[Miw���]�ϛCE�XG�=x�VýK��yc
B^h�j��_��ƿm�$�!.Q�#Z�����z��6�ҍ-��"�~"�b�rE��c�7�ZnN94q%ͣB���B��<W�e
����fh<w�A
�L$K�	��
��~���xZ�U�\��\�:�l\��1��uj���.�H���Y���4�)6���ħ�`�c�O��8��]���/�����X����?��9���˳zvm���=�kV��
�jʫ�z�a�(�h:��;�7�b�g5�ÔD�vN�!�`Y~����5���֛�`�wZe�]NM(9�0د��x�B	W1M�S�q.{�(���%U�Z� �4��*!��C�Lҷ|��u�7*�6�.j�i4�h�����G��(����&O�����q	m�W�C��؇<�&�A�I�������85��r?w�Y�Tp��v2c}�}0q|e�����I�Za%�	��d�����1�X3���Ɖ����T*�ŀ�r�ڥ_5��r����:j��8�[⬖�L߭��sI����{
V�DV�������� ���B�V�A?��n�A1�3�5n���Sp4F�P�&��pxD!�yz=o�E�����k꠩���FK�V77�+!���MF!�~�lws��bܞ�Š'��j�G�����ϯ2�kQ��3�
g�9v�&�c�B����~�����ʭ��^���w����^	�v�~��MV?�2��v4�U�V��ϋʕƗ�����UYT�7T�3�(�%��J�s��]6Q�MW����m߼kN��ks�5ԓ;�-�	f���5��9�$!Ȃ|�!ڴ�IS�o>��G���Z�b6��E�b9���[Ve7n-G&�$��1�M�DT�AԪ�s�Z)��?Xp�5/��DN3`Lqщ�Ò�h�6` %EE�v���lp���6�������n؉���wK)AA���.p!6߳�F�*��z H[�{�S�8wIj2`c�8�ѭ��#->��/�ơr�M+��3��`�D���q52�l,?�h-0�����6P
��<�O� ��Z���O��,	�g �{�^ �18�81�Aw�X�E��rdk^m�Ywګ/'��2fS�7��،�ި�1�
,+��J��O�������2۟&�9 ��|�s=O����ep��zo�E~\���L��(��/ᨸ��K�ƟSL����ʭ�s�­>�%�E�q~q,"��mPnɉ��r���Z�'��3L����`�]y�]����QT�a���s{,��쒭������V'0q��_cla/5�6	��y�]�#g�N��Z���	�M�R)N��bgf �y��pŅۥ$^��7+�ͼ�����y��5���V��xk�_޾fw�	T��?��A�\lt������E��v�q����H{�eC�'�d7[0�֎��ґ<[�/�u�B�/�=�*���Aj��Y�f��)'��?����%v����;DY���Eͯ<�?�%V�aYw���w=����
�܋�l9����Ͳ��T�8�<i�@^Tl��bD����1�]O�i�N~������lL�10Z��9,}��ۯ��X���\q�W���\���SaL�8����ܟ�}G���o H�o��T��y�-%��q��߫؇!�(����=���O�ň��V57n��=VS�@j?;݂�Z��4B6���S�\�u�r�������F��!���0D�t߫�
�"�1nb�BI�K��=�i�� �=�zK2-?�����Rm@���:�u���us�Mx���?�k6��Xn:l�^������|-u�3���w}&��	�Z�>�#zc�\�2e�ֿ)k��0"��^*fNqc�M�d1���Г�>��I����F�adf윿w^h��ߨ]����7����+���}�P�c!������!Z):uC�o��ҽX*�I�[DXҷ���
��ʬ�c�\�LѪ�ʳ�<�o`I���	j��̓j�W��ۥ%�R=���\w��m������}/,�Ѯ��u�ID2�y?�k����Aw;bȨ�=��@�
|���R��w��ǜ�m鼟����O�q6�� 4���{3a�_��5e7o��a?Ѯw1���#]��U��8҇�Ջ�=�d��4�9¿���M�{yy6��So��l��fd����p����pz1�gN��g1\^��ҧ�e�0���n�[���<m5_xcr��87W�%���e�7J���޲e�t�/@�����î�zP�h����*��[UW=���b�I/:T�����f~JŶ�~���YY�^�3m��Dxs���6�H���i�+qh-�;�B�k�+�gWC6t�f�;���0Ǌ��q�"��M��8'M�z&��Ln2��{4L�Ksn,�`35h�%�"��lv��e$~$�4Q�Re9\�j�֛�]CGӝ�9I��/t�����&��-����~�E�B9��r�c}Jc��ΕU�>��rt����G�5��p��������{�j��W��^�
1B1#]1��������-�Q��%�uNF	���f�/W\w4���U������Q���3<��b��EF*��Ӆ�͹Ƹ�LӶ'g�j�=��BEz�Q#�7u�9��o
/��+rI�ްY�Q�[����<�����K��W-���G�B�a�P�hW�9ʪ�������?
�oۥ�߮?�ܪ�ü��Į�Y
m纩���PN9}J}P�V��v1�����6�ZwW�|H2���T�v1q�|y1����Ie�j�!�� �o�����t��P����-�y�(��(����&KKq������z�mV1�
s��~�g��F�$G��LB�c�N�/��lײ�Db�]�k�	b>�&9K��}��\���'o�T�'2(B�aq�R�^}�?���kK���x��ƣ�c�W(��W�#����������=�	@�y��Մcff�urr�����[,�{h�C�xl����C��������(���*]RPŤ�����%��b5�4�r�<v�����+����!��P�/��w/����u����o�@���*}܍Xsp�NH�is�Ҥk�X&q�iޒ�ޒ�o������z��h b.�\�G�0&�}V�#�t��K�"�j!��_/WQ��V��/�b�%~�^�N�4֐W�[�'�ETx�u4��sg�"�(_BãY$)�U�ٌB�%&E��#�W�+4���t�Gb�f]�4Ꙙ�;x�YN9��:��kb��٠�۰�)�����1���9����c���n�CS�1��-�u+�{Ԕ7{����B�Ug��R�X���-�,l�	'�qYf�=~h�<����
fü(�rň>悸mݳ0��?3PM�7맏�T�~��4//�㱘���(4�20=����t��o���Z�����Iz��ұ	Ȇ�]����l�W�^�3���o����b������3�:�eSd��Iy��Ii�"~�p6t�io���샅��2��d%����o��T����G�Ӆ���~_!�Am�a�g���]~�=l�o>����ot�S��4�?R[�";�d��$0�v:��#Z��|;��ùЕ�I�� �QA����I�� }&G�(�ߟ�����!g��T���k"u�kBܻrS�-�)�����
	e�w>YW8����UG��t3���l���3��No��~]ϐ�k�}��N�A�
���Ih~'�Od��iz�Hڧ�S�9�U�k�)�Mm�Qt�^�� �-��U�i�Q|��A/`l�R����6կ�
��F��jT�>�Z�8ҳ�T�Ӌ��e���>��j��֯�a^��l�i�O|�S�]�u����Y���O�
�[t,Vo|���YQS8z���F����BIiE-7|���e��pC��	�G��=����{���C*RjR>�n��a�x�{z�~_d�ĳ�З�H�}�?{��+/b��e���Q΁��~����c�ףI������j�Pe�ͮrn��������᰹�{�Dv����o]�g0��5��9	Yn���v}�]&�5��F��i���2�9j�l	�G���AfaC?�f
�熘�X�/}>�6�Z��F8|���y��Z�F��A����h����j�c��g��3�F�0�fA��{�'���K��432�'�O.�a����(�E�9��Wh���O!����#޽?���:Zy�j�z��)��n��C2Ԣ�4wacq�vav}Y�� �����%��T���:F`�@�S4!$�*�������c���{�Џ0��_W-�1�}���
�C�Q+Ef���Y  ��n�l.�(�y>���6z14��c ~N����l6yQ�\F@Ty�وH����7���X�'��rf�	��e�$H��CKn-B:c͂4�������=ίU�rgн��h��3i�!"�����9�=�%���!�����5�M~@|�����8$`����~{¦4�����~��㿗�j�4Z�~��J�x|������!��2?�_��������L��|�tz;��w��oڼ*� N31����fw�l#$(�aeh3��wKt�$5���с����-��+����v{g�χ�f�v��o��Dl��)������g��ۤ+0�7��hM�$�Ժ�^�?�����$��ͯ6|Sf_�v69/9���m7��xl����r1R�|�|���#Y��Zꄘ��{?�����h��.��aE�Xhn�U�������.w�f!��p��/����:������������c�<D��~xt�k����+\)������|���ٔ@M�2G���t�¾�3�)3_�+qI2���g���-�nm?t�5�*{���<��%饲̋:Ҹ�J�؃*��!�;��"�q7�W�j��`\4/ɜ�K�=�Ւa�(m�7-�zCw��~ ���T$��<i�5k�Z/�@=D�,.���eT=T؂���e��
��,l���S���1F�n���d���_[q@�}��ٰ0�Q��l���_��${�b_1�Z�w����k"�]�^�5�Q��25����Y�}�r��oe��9�������ߩ\���Z�<���z�`ޓEѰ���;��"E�m��5�����/ֲ(���u�gu�V	��I��BÝJ�&�K���>KK�����G����3W��~����8��^�H�`��<u����O�q>��՜D�܄ѹ�/)o�����6*����W����*�=g�/vg]Iw+!-xYyN�v�T�H��0H�5:���)|q.�VK,J�z�������WY����ժ�>�oۈ��^gi4��5��8�l��70�������������	*��ܢ�-1�{���ra��>���c��c��:�L)�g�;�h��w�D��bV�v�הHQe��^�[�d`{�rU�bʊ�:�������+)l����;{�~0�h�zn�l�k���ؙxl��da�l ��~vO���`"��-R�AC�{uƃ�o�3ؕ���~�k�Y������.�r�F���ʠ�rT��D֩ӄӇ�Z�@<٪{*�$���8��AT��a��_-Nos�?���8�q��֮������h�ʉ�����Wa��Ew�r$�Co�T)��sFJ?�`�_-Y�4�b#�7�N��ew���eA��[v������&[/&M��<?�ꮫe/�z�u�9쒌z{QE._+Dr%��w���}��r��Ζ����Û�[$�'=F��Pu��"y������K�F�j��8֏��~��L\�C#����L���XG�������K+Þ��v����|��$�|,�$��OXJꍿL�=l]̐ե��&د��4
��R+��W�����PO���������obb؟�$���Zk�����%��\Y,P���Ʒі�N����*s���F}�m$��F��?�(�́�JH˅<�����N�~�ޯᓾ	���M���{��$�葔,��3�Q��K44]M/�b��T1�Ǵ�oD�AQ!̹7�ţsP��>I�}z}�5$�`$���x�a �x�w?�:ݗ�06e�m����4�i����%>A�p��K����.5�>�o���Z>�hI�+\Y�Q}z�^�<~��D�N.�$�{A���+�� �t(��+����A�<&�7�D��~�'J�5�Ћ�j��a� �K��[���$U`^�Js��̠��=�y�R��E�샱��_*w�����"1K!��u�a���Ó�����_k���U��Hr�u���5e��T��?q�R�:̺�ݰ��C�^�r�b����%�L��Kt�q�@�W��J�Ud�����"�b�;��2�q�w�]'��Y4�މ��Ok��-�g�����
(BD��$�T�H���w�w~�2���p��l`�8Y.1�3a׶u@I��~��{ڻ!�������j��� �\�k�nH8���W��c���>�\�/��0e3��[U�'|�c�%-B*>��=����@au�o��%C1LYp�ϫ�l\������K?�N�1oO�~B���/��է��MK�N��$�bĿ��F/��=��1�R��{����)
s2���s��d�l�,��|$e&̜������{ ��{I2S�ts"1��n^ko����T����B�I���]zv6�Ĕ)i���%L�[�2�i����%��@+�2hҏ���v�h��S��f{h.����H��X���U����G��oR�rTb��ϓ_.A���h>}���N®*���Zp�8��pŃ�G9�RE����#���ϡ���ҏ��TA\�CC�(Ў��~/i����eVf��
|w�#̶��Ę��&�.M�B�"d���Z�|vM�yr3m��4����h[ ����6SaD������y/]�9�0>����g��������;�%Hj/��܉��B�1�G6���1��N�'�%��X�Fq�e��96m�&�E���n j-k��L�/�}�|d?������Z>��b�y��roVqqd���`�T��ғw�p:��U�z��bu%>���R\"N�M_��s�R��eo�v�#�%��㖴���|ί���>-��$d��8��Y>�du8Y�)M�>/);����I"��}a[�zwL�n.L�D��w!˟<�G�ӿ	D����5�|�%��9���m(��mtػ���ó���_��e��g}��	��{G���%��[�w��Z3x���2��m����(%Bu�����sњ�����O�%X�|���N�]��S��|3�������s�?�F�r����3�����N��:E��imB/+s���1r�%�N��t�kG���m��	�����?�����@�%���k�FL���u��������?:��*��)n����;����z�Ht�l���U�\{#��[+���&��'Q�}���4��Թz+k�k!�N�+(��Չ���b�c�7W��mud�?����Uл��q�����@���VRB)i��KRJJ@ZA�[@AI�f��������s]�˙��콟gŽ�{=kϧui���+4�9��^����]	~NNy��|�V�3�H���;��%�]�)��ٞz���+qĽՌ�"ڰ1B#��0e��9�Z>Z�&�1�p��k���|���g	�n �`���Z&H�q����6s�9�����p����$S]�FF	��HˡrR�@�у�	��dB"+��ǩ�111f%�cqSTW��иq����<
����j�:oah"��|�]���򕢭��H�7
F那}�IT��O'6����0�f�f��u�x���DHqΜ�9���|�¿"����ӱ�qp̛����������/�_����<A��Ҷr���mɗ�:k���쬀X�=�X%��k|vS�˔@��$�R���w�qs�k �9����y��dl����^sr���2��d?��՜Ƽ�/�V�6�4��t�B��.}}��J�̛X<��ix�n~�z�/'Q�7`0�d�$�mM�m��;��#oWs�'~�Zp�3�3��x�����x��˩_�[���bZPpUI-;#��@��)���I\1'�����w��[қJ"T"��Le{�r�mkT��el��c<D��`M��'��S�'P8�M%A��<��Vv9סZ��ժ��(r��O�%�Yb��*��-�d��c���F\�X�ӯ�9�k�"]����!b�U���o森���5�;oJUzË0��\��?�G�����f80H�(R��*}�QA�܀���{2�ʑ�E��o���py[k�Q��A�)�]��ⵌ�[Q�^�ME@o�hve�I ������>jnn���ķ����9v�=����iT�z&�g�����0A����|K���bHȖ��h �������q��Q%���l��#�Ǥ#$�S4F���P�鞃���L�|�v:�d�jT֜$��Ea���wC˶-[�ⓓf�i*cŬ���/_��J�Q��t����v�ϙΉ�k�����k�XT��sgx��2��=��E�À^B&"�Z�P.Lr�VZ�����$����>�����^��T�H�j��������;
�QQ��O%���o�n3����
�M�H���;@,��u����z��E��f*	9�r����N��/f�3r����7N��j0���i��[��U�#ߋ��F�Cq�0����4�h�p�32�$���'sG1.H��[_��N=rk:��]���K�忖`6}�5#�XL�ؿ�>���7� �}��#�7�]��<��~���7�^��~�?�áWLzva��D��,�"��������Hm�����׸j�4!��-�v��FjH2��#�Ƨ���|��Պ<�Fs;�q���ʓ��x���gW�Ј��o��K:��)��>n�D)>�gl  ��\,�O�»��+L��|a<R������w���%/{
���H�m3�u���'14��N�V��p�z�.Iђe����IX�;}3;��ɖ֖09�_y���T۳�ɼ�l����O-��u��h1V~��������`�����ߕ�?B�u�`={sN��U�������t�Ē��ڇ!#O;��(K�#
��'M��;���π�]����y}.^�3�g��>C�/�R����)_�ѳ���e��"߷��y�r
ǝ���Y�3��y������*z_�j�%~��8.N GC�r1�3�li�������	�"��8<S�D_�UL��NdX��$	VJ5�c�z1��o�C�a�Y��=��W&n��h���z�lۺ,�}�W��
7��'�O�L/7�z�d��F�J6NNטi
aT�Z1�lY܌�]K��+�����X"��}���ѽwy�gӯ*5=4 ��´�Og��T�Xg��j��<E�:�bD�c�SB�)�*+
\�&�*kk�'LҨ�L,��,�h�c�P*�ȉ]X���'���O��B��/xH�ĦWc+a�嚜�m�:��X!�K�tVͨ'p��x��	f��t�:�WI�p����2Ϩ]A3�Pک��}�̉�<�}fNIP֩^��%:����>�4r-C�nP�3aa��e�n���>�W-]&�}���FEA�8�$����
f��G?���A}y�/����=V�C�ɡ&y���*y��=���#I��X@��_2�2���Y��������sN�ͫŧ�䦬=v
���6v�V����7�3��䁗,x��E7R�m�yڢ_�K¤6��gv�š�>���ޗ�T�Z�Wf���dpŎ���Ytz��PN�!d0�~aB>:��}݇<G�bb[���1dH�r9���ٕ��f��|��c-�N�y�-�K�{KT�7�o��y���c���U*#����<�Z�)�������P�y|Ҩw}�`�˰��H�;�gedyFK�"Y˂���=��f��P�_��zsK��Ȳ���ۍ�r9�%�]���Q4�D��ת�����34�v��{k.��N�����Hۆ~jC���[�����7�p�U8Ŧ�܄X�/��e��+v��k���f��*��%BGa��3snΐ�z���y�_�js�X$Y^����j�����5�b���_�$�!Y *H��O���W��i։�̲$�2�̃ �i/��p4�V+��!�Ԋ�_�%�pB*��(�[j"�]zC�����QF�~�����ϳM��5��<-ojZR��s]�z��ر�g-OH3�Pl�l��e�Q�L�c�}� ��4Qlv�;c�X=�;~��m��B5���&|+���=��o�!K�N�{���J����ãiq����)x��R�Y�"��� /I���gp�>%Sq\�=�a�'�mG!���]dZw��_�~$�7{�G���\L=.��G_{|��u�K>�h��a�fȤ�"{4LLCI�W�p��	ۥR��ڼ��4=)�lV����t߱}տ��i�lp�A��}o����ǄB��:D�K\����H|�8�pPX����E)F��'v��H�Ȅ�3�����lŧ�تZ�R�0b^@��aj��3{�[ټ�Fƣ�^rh������HǼۘ[���3����E+��Q�>`d�����v5oݼ�
��s|�'\����� �Oj����#���ü����ʤ��}��R1�kT�{PԤ�����U>�Lt�.�L���$�~T}2�@Pfj@ �9������ػ<�i����\��G+�������ͮ�nb�I�m��7?�!���X�9��>�W	�oQ�c)��j��	=�'B����zd���_�9���b[��ν]N�[�kp���<�1"d��p�my�rJ�������.�k�|���^\��n���Ͽ��/�������n?���q��˂>�b�mJt��*W�Qj������5ċ(�������Y	��:}*�߇�Ӯ�x4�"pZ�ua\��	ԣ	�O�c�q���$��G
9��ߎ�	�̃{Y���r�@qSݐ��{6�.���uy�;���-O��_EFF<4�"��˄S>����0/��ѹ=_u3-J,?,*��}~%t�s�^)y���u*1����u-X����'[�L��?w�Q��U�W�q�V<r����W�Hlp#5Noۀݧ�����G(3t+r���z�[���o��k����9���>D �"k��}.Cg]�g\J�cj�~ŕdC�Wl�Lv��8��ʗR��YW^!8n���z�/W�p����������n{w��E�Cv���[�m��I?���J9?1�G�rj��`�Rx�vV{^;���K`��C���/04Z�1ܲ/��٩b�j� ܩ�h�F�hM��%f��)�5O/�m�1�U<��^�)��\�J�F"��Qv�+�^(��r��*�̠Wf��]�o��d����\@��i��LP�=����ދ|ݖ�1������M~&f�C�9���#��˗d� ��^� �'؍f.k�q�Ӳ��	B���Ă���̮��;�4��d����>��$s���"���0������O�7���62��	�||�
c��%��W\�!�^��EBN����L.ﻴ��w��¨X���೏Ko����؁��kЏ]���z��M4B[�@�kE��|�%��;+޾��l���P�I��7�o�
���(h��O�Q�Q�D�ÂP-&��j�E�W��R�pL1<����b<��h�~�yt=�Ð9ۊ^�<\s��Y^�*���`�oZh�: Vz��^��G���wH$N��z����2"�N��	P��<~.�`G�̩�H�"�B{�%A�o!��*/jf��?������!ↈ���d��t*�r5�gE���+E�h�#��[IO����9�H���v�@�@J��0A7Ҍ�Gb;�{ ��r?�|���ؾ�2"%4c�2z�]P�C}�qο����Ì���m>Q�DDZ
����M������ZD�c�R��֨Q T�.ג�p@d8���b�Ʒ����,m|,���z�U��q���2� �Y�z�jz����u�U���x~r�ǱHЁ8rK�A���ߥa���E8���%�`@�=HRB�6�(�k�^G�z�����"�1Oѻֻ�;���/p)	]&|½���y�k@��ȗ�E+r�!2%������Y�6Ƃ^3�W�%� �i��W���$!V@���2UK��)��R�F q�K�X�G&"*�'C؍�<�u��6�,�Y�����Ɉ�pQ�`d|F��KQ��RV��1���q��tZ+�V���������'E�JN�S����3"�B�'^�!�1N�����<]b p�]w�X7#|G��w���P��b��b���v�S+A�8�G�D����2E����i���u���Lq�ciQ�z
{�p����^������P�4�"T�������?Ҡ��0�w��w��d�.~�}n��k�D�}Y[3�oj:�y!J���Lt�15�1[�Ds�  &������䔔��Ƿ0���!v8���GQ��6܄es1��ϓ�/��&���q		�+j�#*����"0*��He���pq!��Ձ�sX88���� �U.��:<G�+0Op� �<�ۗ��t�߿�T���6��cA�g��L��.����Py������#��0��� �����c�����-MmǄ�|���(HbA��.�/֞��oxF�L���[W�p}7���P����^DV(����Nd?ʅ�h�F��]&2:�<b'�EJJ�߲	)��X�T!���"�E����(��2��aaYRIkv T|�bT
���pn�ށ����M��`0�.�"�!�H����b��cS�

�� ��A�_x ��#`���&L����h�ɸ�����#����j����e��J�J��[:H����*�NDX�j�!jC������vu���7ǌ`P`$�%m����, 92q�w;bĆYr��S�p`
H �(�b⃙]��z�lA��	�6؀��$� Ȋ��s�Ѱ�YI q�
o�9�e��4����a@/�=տ͢I�&щ.��6R1O�K��rEϼ�ޫ�H�w�Sv���K'}��y>��FD���u���~8�b�E���"����x�^���9��._� s۴�� v~}hR�v��n*�-�l8�MW=�Nݫ��*#�,Ӻ�E2��e-�9����g�Q���	�~��=��k��K A�ؽ��T���U��L����i��$�y��ۀ���S9Dm^j��|،�w��]��+D�꟫�&>ӡo���%,��iu��P��R��	0P5��Yq�(,v�lw� �V2%ˀ#|��.�#�C��	�I,X+�G��` h͡e�O��.%��yfI�~�\�	=WL�41�mf��s����\�� �)�Ҁ�,���W�	��H-�F_=UN�HA#
��1��"}9�9����w���� �%��������D����^#�{��Uk�n�N��� ���d���_>�5�9Fa13��M�D��ɪ��pfu�N��v�R�q�s��G}�E_�`��o�� ��}Mû`T�h�'qz�q��pɨ�R���l��2\B�Y
.z�u�8��g>L[5d\&�Z�*�W������Hɤ�����﫳�F�?�m��Č*N1]���'��˥P� ��Ml�w����q�9�G���+ \�Ф��o���l����R��x'���¸ڢ�F�������w����t��5bxt�{��'U�+���5~3��m�|���V��ۧxA���逊�y�6�P��v��?r\�q�w��"���M������Ja>)0����2P�,�e��2�5�1W3�p
�茅ϲ�f[M��P�`|����hB��o��o��%o��2�$���X-��A��p��n��?�A[d-ۣ=&��;��Q��4��;���`«���[<���Qh xY�ժgf�utp�0�K����c�|$��x������ o�F_]�A��g׭��[wF
΄u	�L�!-�̗&�������xms�&��f��$�ڊCQ���W|T�ɧ�X3M��L����`=*7V_����s��C<�ob*^Ôg3��Y��)��+���K�sg�y�W�����z��	{~g�2QS����{i=�`�($��A�D���C�6���E���<2��%�r�Zq�&��@�g�o��OsnNٕ�6����;�R���)�s�QQVkHs����"��6Mei�M �<��;���E����[�TfTq�?˵XT+��Ys�۽^UQ���2�5�Xƅq��0�>b.�o
�R]d��&���M�'���$�N,cA>��8���h2Q�.T�a9��Y��}�js��ʽlӵK���$:�T�����Rs��hqa	��eSX;����M4��n���B�`��>���:��������u�d��B�2���f^��X2���Xa������9��\�.�=��)��)^&p|2�H��ao?�"�贎+}��m��Zo�`7T�A���[N@�t��LծJ�����O�V�61�=��3}�B�5�r��}����o�ŵ�;��y��<n�QQ�%��('�X�8��l?�u�R W��7����;_�7(�Wd�`��L��`���R�[0��.u=�}�Si�Q.�{��<Rl���L���kX�QP�pU�dP�cc��~��M�6ҹ��%b������(����Oqf�&w�6�[���|4��S��e��eM�� �PU �x���n�2!��R>�Ｔ�� }��
��~N�z����J�;Y�H�yw�����=�<��j�\V�.t]\������|���=�UN2���h5����?����D���k{VxS���u���E���i��,J�4'vt�ޖ����|�Cj��a7�Qf��#��F��8� ��U]��<��l7n�u�G+�L �(���/*��zD�C3�%��x4CO�o��q7�k`����.��X��ZDz�R�U{���l�'�����&���'�ċ����Z��5���n�mg�m��[���h]x��1��G_ώ^�O8B�~e��I
��m �\_jF��w*��8��5�Ĺϒ����/�qz.Z���چ�	ϳ�@��K�z~�D�x7#�Mӣe�>�K"S�7��b,�i+!�Jf���R7�ԟu�\������
qp,OLG��8����1�ڑk�0��T��L<���!�sR����Ɣgc�<ݾ+�ڽ������J�Qd3��X���w~͉c�!]�+�6��_`t}ɹ�������v=	���|�^z�y{]���wP�b�G�T��a =��}��(N�u}j�2�|d���w��n��ٱ�����w�i���O�׸ULk|�N�Ƈ�h�󇘉�L�P~�$�j]K�8oy!}�����o��؅����W��oݟ���*W�����MS�/IL��0��$f������:T�p�%�����?���z�#�F[��.@�F��I:[���8�3��7�]h�%�!>�
PA��T+T�z���/`�$>�M�Hj������U��58ڡ"����p�/^��|,�U��᫣cݴ�w|�U�JB%	�����LM_�*V;����#qa>/�R��u��N��M�FO��J9ˊ�j�?���jC�*�����|Z�8Ύb�i�����V8k� ��������$�C'0Ö�o}�r"c�h���:�'.^�����K�9���f�9�ē��C�y��ؚ�XӇ� ):E�5(l��I�IIDq��A�y����́�inr�?r�K���8A2�ԑ�;a����AL�B��]�E�Z/_���հ�?��r��c��<g���^y� "M/2cjX�t��C���I�N�����}b��ř|�@�1Ph���d������!ԁv4I���7�����D)d�;����CHpY?�hޔ��/�`��8���q�9.�38�R��kg��y����-��O�=�;|\�@��D��;X_�D��	w����Is�!?� ���a���g���^ݳ�<�Z��Y�h���~YQm����B�{[���/Q���+�8�XJ"���GZFJ/'ޅ�
��1�~���b�w��`s���]�a�b�fW������is,,6!6.ސ���ٚ�3b�'ʏ����\��	GNLhzw�������EEM�o֍?4;`�R����%6���kk���{�x����W����wԿ�����#��o��m��%�<U|X���- �;c�{,����2%�5�;&ߛ�'���f8qej�������"~��������\@������Ջ���X��\��yWP�G�ɵ�GkR��w�+�M(/Y.$<V�W����Y���w��.�D~]��lN�����l�pܺl���"��>�}��%!Ԧ߇����$/_�s�����5�$}�7K�N;vp����K?��E:Qu�������6ϭ��������a�lqK%�3Y3=5�b=(�� &��Ӊ�E��K����Y�	��K4̿�����/�J���j��C�aO/}���w�uwwOʆ\����@����m���o��.v�2U���ede��c�u���)��=��Boȕ��!��m��iI������Zɝ]
��z�xn�7�#�_�ύ�DQ+���1��w�;�I5�|Z����4�v����D�V_��� ��(�N#�!���c��)�D;�pg�wq��q��TA�.B�F����)&��&i�zв���(�?#����Q���kB/�ͣ+�2�=u�o���s]�ty�>��}u��|{�V�A���f�+�W8{
W��w��Em�;�o��a�F��O��=��BKT�
��7U[���#����?�Kҧ���a7//P���Ȫ4چ���i;#��;�lR���^y�DS��}�s�q�)��ٮg6V]�繩�'tc�;����3M��|ְځ��\[4'$�)�o<�w��G�Hm�#��T{��"%���K��s�:l*�5o7H��M��L�����>�7S��0U?_��/ԏ�!�	Cs����Bs�-m-5-U���>*���Dz���O$P� �뼎)�E�/	F��y�FO˛0ATꥠʵ��G���s�
S���$�s�,=ok�&e���D_@0��#k/h����j�e��5K�Nj�N�����q���bc*kqٛ�eU���$�*���c�r6���? �_����;n���x�Ӝ<�:���g�:/�t4��T��[Q8JÐZ�a�K���3֙�$�Wհv��n���ǵ�˯^�����o㉶��)�w�T�}�t<�_�.�l#��C�r�R^-�iǐ�4��W���
��ʰ�k�$��3�.�ۘu��ji��Ox���[�0�4�$�^w0Y�deQNOO�{D�$�{iOth+VrҞ�.����r7�M�h�sG���x��*���ʫ���f$?�k΂��Թ��5H���t�x�C�ܯ"jWb��q������ϰ���1��� ��+*��e��U ��$�Z���J�L
�����[U;]�%�(Y����<uڧ��,x��d�'w��i-�ϫv���?*�Y҈Z�e��t��,����m�m?(G��/U�������쮍m�E��h�)�������e����� &�&�܋!�F���ɗ{cФ�}9��`ʲ�!�K��%����we�SaҬ%ʸTH�s���ʐ��?ò��%��a1�1u9�)5�_y�7�UaNz�|!��O\!��� �A��N��E7ڇ0��9V�l;�o���i�}O+`�ޯ�ji@�ʶG�\�NB�})�u���8���QmȲ�3Ϫ���Vl%�K�e>�_֞f���G�{)bE���gG4L�	��'h&9��Y�O^���3HBu6F[�Le0�k��,�$?LPݦ�1f*)F���IM��$%p�I���|beL:��m�o`��������~��\�(ƨ��<]A�ns�2"�(��34}��F��<~JF�����cRh3#�����rQ��|L,L�8���|��W��r�ڹ�G�0�3�O�缋��c��폈�s��ڀ0�cX/��q:k}صq��<��=��������k��m�v�x��Ş	)lo�p�A69�,}���p�B�hl��ԗ�6`.��|u���*;��Nq[�\\����g��ψB;0_��vDg����V� ���w.z��:&�|w篣���o����:y�V��'TE��9������B�'���O�ޮ�,����[i�vb^P�t�>���u�.ѭ��N7�C�ڸ{�V�&�5X�/nw����g���e��~w����)��z��y£����s��8�Iڬ���*�h�,+�?'����xswJ�!����Q�����r>*��w|�e"��:%����_��9ָ����3yu�h�J�&��'�Ƙ��� n�*�}]u�!�c�+��B�u�f�����5R"&�E��Z������u�ŋ��m�d��?��+4�7kb��>l�{U�E@���Z����<�*�	�!��m��2���v�2�S��J;U#�g��P����W����t?�\)	��N��i�»��)p�f6�/�.���'DIN��]�''�6Q�"vL�䶓�vg�K�y���Ko�����ڮ=˰�՗��m�ٓS��[PI!����ƫ��¨�%�:pq����=r"�uB�A�U��nj��D���;�K�ڸ�&�`���)"pe6�U9����5&'����G��?��6aM(�MF+j�ż�_ w�<�b���""���� �!tN�N��pJ�9�T�vF�9��rTq���﹉��聛`�J��`EK�,|z��A���vc�4��8��'0��XK��_�@w@��t���da���F��jv��O� ���v^	�1%�<͍��,}1���1֎�N���h�H��z�j)���^���垭�̿8`�|W۱qW (�=����V�Ŧ)��d��NN�}*Y[e"��x�?o3g�.�L��sT酢9�\Mܮ�u�$��nN�D�g�L��Z*�D)A5[p�#꼈q���|�4 �/N
�����|z)�&ݟ����L4�X��r{hB�ĺl?	n�xy�@�&͠������R���A?����K�Wg���X��V
ِ��g�3��]�	�µA媨�(�����T���#��=�Aci��;ڥo��ɏ^W�!N��w��IE�E��:7��\�9o&k���R�]�xe��:��gg�ҥU$�PڳW��0���J�ҏ��x�d�o�������m.H9�Xh�gY?�	�V�������oc����
�.��_����r��)@�2� /���2�<AAH5���",Ѓʗ��P�[IH^~�H-����[�o+�~2]p΃$'樂�+Mw~�]�c�8�m����$ov�+7��|D[?�wfoj��m��˨c���閍g��	� L����f�v��q�f��Y�5���;l9�����)9�s@ۂ��#��7�b�mǽ�E�`�{ꧥ�7 ���D��$Lqx~zn��ٗ�o�b�U�W�/]���<W	�8/�U��'$����c��9H�z%����#(��yM�9hZ�p��{�yָ��w#�Gj�'U5�?���⢏�Y�^H��h�;;���Z�̎����S����r���䐘������]���z�\��+�/5�^�t1��8LR �[-S,�lBЄ 'U��u���ď�W��R2+K�{2�6W�8�#ve�Y��D#IȌU�hr:$Dq��^مzW���%�v8Q��Iۜo���o3�w�Ȣ�E�m�A��j������&o(�?Q�[���{{�g#�R��7�����߱�����F~4�͈<m�0 9+>]�z,%�Ξ]�^�"S��py4���E;�!!�Q�'ٮ1I񽔫$���s�K	
���A��yU�x��B��4ψL>\���1@R�6�UF���P��4tnCZ���b�M?QKS�MU�R�cG'��c����03/Z��HK�t:c=1��̼��a�f�nB���"�7��3�⼕�rS���[���וV����bfT����Mä�˫��!�Gj�y��ο���eZ8��9���ޔ��4��ͰpĻ�������Y��X�0����ٿ*��F
�I(��ߥlhV�u�͊�*1���lt֦}�q ��K�%F�	O�K�i��P,wLG�*�L�T�H�/��8vxDl��e��P���A`k��C�wը��7�@��@��dKJa�]�ij��.۽�(��ͫ__��?p��.�e�z�v�޿�Y���?X�7+�R�G�
�#�R��s��gVo�Q����՟�(��s5�g��>��(RL��B��v�Σ�;rp-)�%��r��(��3�|����xO`��J�[�~Ĺ5ax,H��ݛ4���V���]d��RG�:��k*�Ỵ�bC�~��ǧF����K�%�2���Q�/.�CU�Y��xh��q#A���P��]ㅴ���U����`k�������cϚ��s��'���t�G����iD!Nw������t%�F��?L��y���1��b؃n{NLU�r��K�v҂�J�ܱc/����Ώ��
���<��*�i�d�U���~j<.M�����wW��:Ї�a����V�Yb��`J���3��(`z��ԉ�͢�ȣ��2{�cq�fN�G(�{�����sS������(OHڢV�0���)%�P�C�ax��i�Hv]�(��!� ni\�f�$���*K��\��7r�E6ф��σ�B��@��Pɏߖ�*x3y��W{�>P��-�0C'X�H2\mo�z��9:�t:!H�e��5�q����k��3-�>O�z<��A�Ӯ�:���Q��:��Оyq�i��1�xH�~���O������!m��o�����ֆ�@����*�)��	���C��
n&V7��L���)��
>4�^�y�0s$�ǳҔw�]�̭}5(���"���h s���!���xjǣ�y�=��g<B��Ǡ��9P\?7hX�l���j�#�2�캹�!��{�#g)��a�:�`zFs��Z3�����Zn
��:~����k��bU��ߨw�գ~8�S��m��{�S.&����z�s�����������n���UfkuĪi)s� z�Z)J-剼�v0i��Zdg�~�� �4�zp������a�d
{I����k9uU[��Í�[&�oL�V�=�VhX��� ó��JV4#H�
ў�����Y� t��'s+�d�g˸�J���
��}�;C�J��X�M�`A5������2ʾӱ҇2��RN�<���+��/��u�vr񭫆k������ٟʽMh�ؾ׀�%m�jV��_�^����rUն�ܱb>`'���0O�mS������!���'^������z�b1��Q����Xx�����l�� ��[H�:>��Q��4�L�ti1��A��g��~I�7]�����.[�@翩3�Zi�����'f�Jũ�4)�]1,��卻<�k��+[�BS�j)B������\>G@�w,�Iџl��j��r��N�$M�C�X5!�m�tA/�BAs,��0�B�}���ǅ�I���M���?��E������N7��ĠRIkz&�¤����_*t���iv)H���Z��a�耭6ޝ���<>	�M�+��Z5�*��eǳ���O~z��R�Q��4qL�U�����|Es�qI}3N�D�����1#x��o�e��RN���5��s1�,�^�,���Bȕ�������lNt)q%=����'?����!�M�4�=	���E;��`�L4�c�=����R qfW�;�� 11������$||#$�{�?��&w&<�rJ������\?~�ݒߡ�\Kܟ����&<�0_",�#���\ka��"��Z�q�;y�[0Z%Q��oϻ�=�\��ؼ��5���Ig�Y��[t�
2�
PXQh��k�(���Պ��=qi��7��6�>sn����a�|� ��;[@jB�z:�U0���`����s�UpP�G��a��TK-�0鋕"��=���&&E�y�;s��i��5��gx�G��1K�����s������5�L�O��v~�ku5��!9��
[��&��:;�~���ڷ��R��o�ᾯ��oa��S�_ss��~��>4H��2����Ǆ��R�[C�~�kQ�^yt�o#,2�%�'4[�@Dь���H��ո��.��Ut�\v�l�	�e��T�6APs5��`<�l�O^��a�&��hH۾����^�b�^fꛗ�=D��M������9ynǌ0�	�W\Ml^M���y8Q!�~*v�[U�v��:�s�t�@u8��[6���;-�=���jj���$�P%���K���;�9
	
���D(W��%+*t	Ⱥ��x
�_��y	bS/a�;�]�$����zh�(�]��d^�(�.sXD�57���M�a~����J��XVG#-����/��*����⢋P�������&S�M�A�i�\���Sl���H�ʧԚp�l]����_��Ƕ���4ԎO�����:���d�]6�^1Cfx0ɡ�p{]O_y���U�t�|�EY�X�[{P�&��З��uTZ�R��k��.��p�m��>"�V��e�kr�y�����O����W��H������I6���:>:���K�OXx=��K#�l�?��.���
3 H�9�Ԛ�:�;�,V��u��$��>[��	I��J��"~_��]�,��♻,��n���&mF�b�S�W��ʡP�<-&6�|��p�����5�r1[�^�V���1v;��G�c���b�����`{��?�i���a���D>bY�\ey�9ޝ�!L|x
ߣb����
)�[�����K��ʩI-Ϫ�%� �� R�\F ��61�����ar��$���< -r�����{�dʊ&[�BPnj!ǅ���5e?2��!K��8M6�?�'<�	��}�F�"�w�����n�N�ځW�^���M�f�>u�����Zmj��v�d���j�Y c�W��!�WL7��N�P6)x%V��0�f��S;�G�#�[����%4�����r�a�3���^$�����!DŜ����
��0�$�s�m�mƏ���b����o�?��V�*�9a�p���c
��<����"�*D&�A��D5�-Tcw7�;�I�����d8/+M�=j��T�}n'���eO3C~R������~�B��R��rlw3�;��u_�U����<Ϗ��IB�$�{���f�[�o�f>j��|���u��68��ꋘ�E�A���� ��&<�8��B�Ll��h���ѐ��ؐ�;��n�袞Ue�c}�
��!ʻ���� �"�k�<���'�7�K���H�6p�М��P�H>&O��(�N./;z`"� �F/X��F;�����_^^*�����w�j�:]6�,�$�9�Ζ�|,�?��@3$`�$�������1W�.��������4�J5��t���5�Ƭ��8p�Xf�N����;�MC�������>�7qq�W�~�o�Q74�� �p(3CUFg�p}�$�7��NH�_ �>v�F�$$�0�;��&���3{�
+������V�&��?�x��B�ڊI~�q��Xnb�\f
�pO�t���Ms���=��]���k.�-zp�B�l��3�Z�+4��5ʒ���v�Yu�j��c u���l�{���wƛ���تb�Z�XӍ\o+KS	�ղ�
!���;1�$O;iC#�Y߉�
�KD%���0��l�wvT,j#�����V@U��4�g��}�����ؓ�O�Iz���:�G���� 6do"]��;�ܷ0\�7�Y<I�Ĝx.[{��-�ȠJ��Q�d,֔w���d|0�޷i8v�k�*3�o6�+��f�;~LQ�g��B�[���k�G���t�3
��i�0�ֿ˯ЎUnj�G
WHH���C�ٹj�8w)~��0���㱇�zh�dv��EUP��Ȋ{�z{X[#��u���t���w��xd�.E
w #�L��"+Y�l��a}�,���	X����f����"G���K��H�>I([GIP�C���C��
 L>�4������Q�_��WR���<@�6�Y�j����u�g�����Tpj�B��<3���J\2���zS3�c�K�s���޾��!�����;�-$��d{yK�o�X�����������&W��d@ŹUhm���&�b�bke��p���s6 �a5�ؖe2�����)��	�ݝ�$�5��Np�E� x x� ���.!�a��gaq��[����Wu���E���3�3��<===zW!B{�� ���@��|O�K�]�*Hۙ��j��m��5@�F�E�bj[`���S��y�p|�(m�m}��$Mno�"ձn��D��Q�1���H��
6O�ɭ�N�N�*h���jF(1JA��H�wB̻�S8tI�ˑd�X���e�U�<a�.N�7oQe%G��.ڛY�-71`r�������R;���#��8�{�|zCy&���}և�Փ]$�Ȟ۽���5\��Ue�G�8�0@�1��(ʠ�
D]�c{����}6�Y���MC�嫙*q,k��&�yo�o�x��΍ٽ�J�6<n4ݡ�RgA��(p,b~�M-
����4'�2�����[�|�������:h
�	�e�����{"�S�j䉚!"^����Ə���xk�k��f����qyT�xtsW�z�5���o������&Ͻ������y^{�u�2������?z�l�W0J��^Z��wz��n/	h?��I��Ҡ?�ҙ��L��,��mS�󠴬iB�y��������a�S�7��
S�}�d�һ��7��}���.��9�'=�v���4����G+�r{�TJ�MK&\W��.rb���Bb***-��x���� :/:ȼLB������
N'6+ ��V/�-/X�n!��W��G�
3��Jv�j�4陳����[��G:�r�߽bC՛�6����(1�V�T�����}�ήn [���e�(l>C���
�V��JTX��d����\��}�o%
�1_����[�F�F�-�%pt`he��^�^QF�Ł[�u��s2u�{���;�aP�oBU躽I�v���N���+�K�|��tq~Nf��?�US[�3w��P'/((>q������	���U�Od�B�9�v��QsT�>w��$��n��y�wU�4!��f����d͝�T����~?��cp:�'j�¹��.3c����Ԕ{�y�'id����l=Ëh�숳TG]p1D
��ǌ���%��"�Q��"�W,���;[c?*dp�O};"$�V���i��& 3�(�z4� ��^!N�vŏ1?�������|fjj���n���s�lM3�Ӣ��O�p	�f�DP���)����P��߳���`�v��o�:����!Pgؠ��X  S�24�x�ď�w�h$q��ɗ�����;7vxB�/<�����D0|��-(k>{({�-M1�}Y��T��?�X�P �!xr�� �:cw�Ai�Ѭ��{����lSY�[�|]t��^�y9���ȭCn��P���#��H��·b(N̲�]á A�z^c'G!��G�'*�Co�e�mr�e"y?�>E�YL��.�u�4vx�L!rq@T��rGι�`	VJ�+��� ��]�����U(��ĩқ)����C|��I�/q)�����ʭ��(�zi�)����X_�oJr*�������]�YuAË�끤������Z�ϒx40jݠ�P��Æ��56�X-_Sx�<0���r��aT����v9bȐ"�-#��Ы'y(5;Bb�}�ϠH0�s�����y5�}�8�-��9U$9�F�\��Mt�1ަ�i��V�rQ�W�=𯏄h(��ڞd��'p^�O��.%#_aI��ۈ�{�Jb�G��=��Q��x��Re�h�k��d>?U���[��{(�[�
�*)�LM^���c����ضsS:~u;�^�#Q�8�aO��_M-{�H��ӼRqG�z�{s�VY��1�x{s`	?q���.̝Q7�޳�ɂ�#Ǻy�Y��6���h6���	����=�ٜ�%���}W9V��V��T�`t�RSn�����o�϶.Mo�{k�ȍ9I3Os`h�/p�Ӄ�A��=���j j���[�MdZ���e�m|����B,m p�o����_�~�$��U�G(��>�#�u�6D{��9N��~�o`�G_j���Yuɹ���nm\;�o>�¶��Fn6sfG��%܂��-1V%ê�������Ґ�U��N��,���+ġ#?s���=�R�U��g�_�(tn�$tA�;�誼��Dl���i,���y%"�rn�%H����޽_�_�j�:Ծ:�TAf�����Dh1��7�H���2D�t׌Ja:D����o�1��e�W��5�"��|���N��:���g�R�URZu�������|9��"%�i������O���D��0�4w�R*�S�5�3�C^{��i6��j����v�h�^/��	is���ڐ̚��1���a�MR�U��N%wOE?][l�>��RW�)��2tC�|-ƲdG���f��K�x�!�uͅ���'D�p�� ���krӟ1�n�L;_��ܺK7��o*�?ŝ����Q�O�j��>-:ZT�7[�r�jƶpX�VT�|'q�y�{�^C�r�Zr�(�%��)�R�({�ĸ}���O�?*7V)0/Oy}u�}�	*�zS^�J��ya5���Sgi�ܱ��*��OYԼ���7��l%R̵S;��9͂?�;ޞ��y�/�%����t�ָ��bG#���{c�?R���,�.���9�R7�!���5�!�΢����-+������m`�cn*'���ݨ�В��5��;��C��+֛�?�[ Z/��F��W�G}����'d	��t��P��^�����uO��r������	ؤ0��
�r�2�1��SŴ��7-�Tbb}��+u���s�*=�~7�ň~w���G����a�\� j�F�(	d��Qg��7�����&F{g��*�5I�������j�ĽZ:�kr��4UuR匥����e�!�ē��˃0WGD��X*���2��m�'��#x=OuLI��d�dI0恦���h�2����cOl�~��~��+w�<K�(�fȗ�a��4"�!+"�w@���G��EJң�־�4�/�ڸpK7��cT	�F��_�A��VqT=�k�[�O��F�K���~��=��8p����_�b��T�����2Ƒ������D�����с�SE�����]���x�Bl���� f@f���Q����ʫa����/��7�!|�?X*�$�F� ?Pzv���d�58�B2��Y3��k�R�|��t�\x2k�Ț�*cQ�҉�_�>%�n�������QH��Hy�n�gh%�.IbjsL��S��7��p��F��Q������th��G��`��j2�o��_;M7<:F��.F�24!���F�"�v�V�
��*_��/������)GҌ�m���Ƚe�-�0.���W�x�W�� G�p�N�����Jqp��=�do���'E�m�0��N�k�.�"컊��]��C�������@���`q`����,�d���@�������O(�hDt�� ��\z��f�c�Fn7Dt%�}��Uy�A��"e��,!xc���u��{�'��!�~������l���������{�"6r�[3 �h��`�x\C���C��n����*���?����"z-�T�ƛ{��~����9PV�Ջ)s�J&q��Ƀ�+q�|����)��� H;�ŝ�{n��]}�QE�m0���ƟR�����^���$�4�*��	ND��8l�ҩ~�)��5_*V���_Ϲ��OB�c�ϼGm@%�%N���no���BUQ��-&�C+��1p	6�|�<+'��nX���0�����R��L����g��-�w��!�>��1�>9�
����!�j��sV�hc�&L-�C�3�wT�H������KG	��|E�k���s��=O'w�y~��{��Kߔt�g$O�/�-�@~�0�{,7�;����8�4��Q.��`��~�����wg�X��H7Mt���k�.���)?
fv/Z![o���Ybt�hT!�د ��[M]����"�=m��O�5�ǒ�3\��)t��M�u2AjI'�&���*j~��^2@��7s�������-��@r�%d%�8��A:�+��_)¿W�r�o�x=��q��՗��T����q��1vќh���5Z����.�����Jě�1���E���W�a\P\�JB*�>s�#��-�-5
3CC��)@/Ќym�E���7)Ɍ9�i��GE.+$D��S����V0񧸷Hlu+	�'Pv%B	���b���
&a�<A�H;<��U��=�F�q`0���� e��Y�,y�1~��7*j�h�'X-�8d��jh���H�a�ˬ�n*8�d�����H�PQ�a[��4ؠ.tn���JCtP�g������|yЙ�i_rb��j���(zV��L����#��t��n^g&��&��/�|␡���1]�jv�8~�������Vr���52�O���yTG+~7��m��GyB���֑�#�(8�&�ڏ����1�D��o�V�79�/����>�������G+��A*B�O)Y@+���??������w-P^����0�%iF��u�~���Cl���D�4҃�W�G�Gs��y��s�3����5�4&o�G,�;8"CO�Ʒ�ӈ0~6ّ>'S�w�tE�˸jA���V�f�ق�����4V��(�n;/��p�!p�͚�Q����9���xx �~k89�����|f9r�W�/E*��)��ѡ ۚDQ|Q[`�-0
	�=���7�[��I�Y��‷��	�'��s��x(�̞F�4�//2:^�F���Rn#��e����b�
��H|�L7�����6����}Xd�l�Q���&����3NuS^����`4}��R�h��Zdyj1֢ʗۼ�%Ў��Gw�����E*�i`k�>����gy�\\%��ud�|������=��{jǛ��a����Ĵ��s���Ҿ�H���<�B��Z��u���z�`h�9n���M^7;2P���s�����= 97�@2��t����҄S8,�u��|:�!R��i_�_<�d���gcC��+�ҭ^�|z�n�)>�Z��4�^*E#�� ��`�V�_�B��M�!���K<�o��+�k�$�y��L/�,��O2}u=%S$��yH%�T�w��v ��Bk�%�,o__
ӟe=ݹ1��������:ɘ��6���(/��3��̃������j�8cq�z�	���g	����>�3Z^���/��-	0�4
�^���o�׀�?t���ui(��%���Bt�X�<0l%��'�}ޭ=���2�3�ijP�Z��}���c��z�u�����t�=��u��T$`G��E]��{	R��Y+E��`K$������O��a�quo�n:󭕧 ��yq�;IJ��f�$k&��9���q�̧Up<�2�$�I�d�rш[��b�G��mU��F�S�("Y���p����T/��g��˨<�C�F�`�E�`DQ	��Hƪ%@ o��[./QA2{�$�`�N�
�c��'����Ome[���vTί�(L���]f�5�=�ت�����Ǉ���3:&f���,���`V���ȧ��w���~i����(��O�(R�����u�䎳��?�2^$���	�m��?���#1῍5Bg{�t"�K#]@4뤮9��%��L�K�3�����#!k�N
�a�$��EpAx��2$�S�O��En�����~��Z&�����#Qx��:�ף띹Ij�\0n���Ƽo���� ۚ��70TW����QGLT��v��X+�tS�d�uc�>/ޭ������Q ���g�82�׷�L�!K�H�Ah�X�|kr`9?���	����B�hpD;5���i >ft����[<om��W�u2v)�bxs0a�|�q����&��O�����&p��H!$D!�9�����$F��iz�Lɻ��OrE�q+Ý�)�ÄB��$�ع�[g舾��c[/��	���()y�ģ�gvM�X[��mD��q��
鉈�_�2S�����?7%��3��E}�T}(�@?22����w����K�H_J
��u���v�SYy����7���U�xb���'/&�'+�V�-����x��� F�<�𗌱��c9�ȋXb�]��P8b�$�X�f��4VM'/��.�a�S���������O/L����}W`�DRZ���xzĐ��v��#�X�V�͒�c����Q[�ˣUW/֢0Z���	�O����^�d�}1>N�k��8�Y��ďY���L���ߢ�^�>e/����v���Fi3�p��@6]�h���*&�d!�����"qae���i|u����JԲ���e^�x���k���)qԜ~!AjY�5��B��ö~����JS�Ym�����EOo�U����(���de����B:Y��0d����G�t2&CS[��Sw�z �+�e6�xYK�6wr����ĳ��l���.�DVP����PK����ho��-���mf��U��E���]j�6����D����g��&��g�WTD �	r=9C��H�P�֎�b�T�b�ږ&&����PL?�������
�8�&��t�$���טz��t?����N�F�[唕u��ɛ�#NE��3�ȧ���<[%��s@�'�a���%-r�AKy�7�?�����N���p�9��ﷷN���0
[��*�?@,��YCFC�|�3��h^X'��宴��VDi�
�7�?m�� �5�8Q���n�����<w(��ey~%�ꋊ�N7�B���oX��1���y'�eK5���py�����55��ݚ��П�8`�@��K��:9D�e�[������v=�K�>g[�l�'��ʚpd<%�b����1b����G��JR�^�6l�w��`	����oq\���O��=���J�?p+�����T��%[�VJ�_��];��|�/��_�Tx[��1��5GXk�?��RFc7G»Z�xxd�J���.8��Ysr���G�>9���ǉ��
�`eo�*��߇�ckh�$*���4��C�B��F�Ȁ���~�+��l�� \�w���Ej�/���01�`��nNB���rAC��9NNVN�;x���|�F�>���R7Gc.ۛ���T�r��ѻ0't؍��PŰ�09�s�2eҺٺx��^4���P����3f�5⎦r>2�yK�8���c���e�B/.@G�ּc�ڧEv����.v%�#�Ɂ����_��F�ʑ3@����H���_��N��p��Е�0ڋ�T�ռ�,�����a$���D�K�����8�I��*�O{������~��u'��i���/j]BD�9^o�td0���w�>��i���,���Sڶ�/���q���p�nd��_�ԣ�|a�C|B�%�f�u�Р6~�&��9�}�\�I�h�wn�$EÊ��,��y�06�A�)蟉�~�m��~�V��J��%���@ք~�`'��M?�+���j�%�*�W��O�a�f��[���m\���`�ּ��}J��@2ُ�P��6��y�M����Eޯ�x���#.
~��^SQ�&�=i~Bڰ�������Xm��?�H8��*��JÏk?f�g����������@�l �Uiқ�B�{v��^N��tu�km�@ϴ�n6�>m/�a�&��+�ǡq�"��?��f�o��1�f1�E���U��h�6���}��5�Oz����.�N�j9aD�!��D$s˶Q�o0�o���hr�S��Wdk���y���ڞ���ό��-�j˚&���)c�@�;����dJ�=�םZ['�0�׆����iw�ͳ/�Y�j��t���{���`k�@b�dt�"漻�4�Ysk�;��q�p&\�&��Q�>��������j���b+P�A�VU`+
D+���r��V��{�n������Ļ<��4�v��~_qκ�\8�1;5�<�������$>>/j����$�?Fn^��X�2��m~��S��r��6�S�9��j���rs 4D5b�"�O�/�֦���댽�-Y���Fyc�/���}��x�	���Q�����6us��]��S��E"y�gA�xrDc�|Ÿ�&5o�V���n�v��R�.͘�Q}~[����נ�A�T�q��j:�[�Ԯ���t�L�`ڎ���&�[|��Y�A���ł�y'�ǳi`� �m�̓�rL*�<�-A}�Lӧx��N��7����}M��b:p��6���ƆB��}�P΄M���K(�N�!����p�֩4I6%�̆
/�E�F:<�'���Tl�I�@����n��]�.��/�z��m5-�n&~o߁��D}����6>����'h~rnc���S�H�Qws�D���w��-�7X��:J"���~Q�AJ�̵��u�_o�h���Qr����>B<����H���R>�p��Ί��ٿ��rMb�[�+bQ���� ۊ讑_e�&���6������3�W�@���w徹�uEٕb��	M�Ei�>wi�$���?�2�6pSi+��}��Z����`:q��8�ӧ��.)$�%9^2��k�(����`U�gZ烇��q7;�,�+�|(���d"TU���7���f)��-t	�:S���y��:0��eJ|a/�f��de�ܩ�T��M\�%d� ��Q\{�n��V�����$m"h'��܆y�Q��VSrCW�v�����xG�.x��<S7�̒k� $H�<�Pb���P;���q<���S�r�^�S�F�*f��v��{YEȋ��(���˦�U�-���8�~kF�.�|;̶NƋ�P���E���ϝdUQ-7L��Y���&���⊃Q�/���G?jmF�+�:����|�лuУg��Y����ܴc�H&R��O#f��v���kԬn��h�
v4�K8
�!&x�i��\W�W	^�9u]w\h�O���'��qg;;oS����sB�&�f(Ʈ� ��J2��?�n�.���v�:���g�f����y�U�����A��;�7x|!�C�6/d�OC1;�E����X��x��E2t�-Qr5�l��P3n?ۣ�6Lz4�hC+�=�J"U�(!�l!��c�Hi���~��L?�-���v^���\�'y=��f�d-�ZK=f#J��� �Qj�[M�3	�:��]݋}�k���g MZ+<�m�Sm_"�@ū��d�l 3)��/^���!d���\k�$>Z	���� �8��fՇ��ٽ|�\�Ӱ�H`����Cy=_�^�T������ͻ���A���ѷ�@��!��|ncw�N"��.;�[3�V����G�>T��5P[�-����,J�a�ƈ�^�`Yl1#�|�x��?��M<�=��;��f���n҃��l+���=��ެ���j�R��缿�3�ъ ,`�ξ�.�۾;@2�e���و'�aD-a�Ng����&7�Y���_W$s=�zp��,t��� ݹ�HZ�����Sp���X~����J �+K��z�
r��Ⱥhd~�L�Q�W�<�]�,`�������6G����`��؈E�
������[�q��ƛk�z�h�I@��	�щd�s��tVQ�V�3��3kN���ӻa8�Ì�� !�T���� �*$7�Z)M��,5-�dƜ�s��\N��ώ�.��y��\i�u|��u|�mY���$�1�R���yQFÑ]W�i/t�@�x�N��5&6�8�?�����#�^�o�������⡮���omMǚԌk��,�r�zu�o���('L�\0��s�4�E�j=�e}7U#d��1�*Y>f�$��@,U2G��iA"�Sќ�#����=մ�-��s�<6^���>��@�cz�WAY�r���4Uu��Gs/I�-<Y��vV#~���yg��ļ���³��n �����bw(#�5.�J$�(�3�!"(M�aD�	m�j{_�u��_��=����Z�����y���d<������������2�{S��a�i�ˎ�[\��6��{R_����p��׿�q$����U%ɗ_:��a�nۜ�Ib,�l]�\`C>-:�غ�&�5�l� f����s;3���ck.%�CHp�@D)R=������e5���	q>�9�̎3�r!w%!Ȑ�$�C3O���q$��|�YClSufy�J��1"��n�9�t߭I�Y����>ve�y���u$L��Hn
�?iM^�xêj��Ez�����>ٞ��r�e�nۜ�L�`;��r��Ò��z^�q@����������7�"J�#f�̀iF�D�c����z�0��ӿd���y͝l�&v�RG魀���i�VG�� H�a��a��qh�0|g���ޱ�IY3�&WC�OF�:����r��R ϻ��wG�i��~�J2���A��tZyBN�
X��aTROg"CO3�c7�Wk<�(.��e4�:�c/�0��a�	M0���c˾��U��Uw����wH�������Q�R\/���h���:}���W���AW�����eS7���;x��cO�\������@�]q�$�Ski�uKaө�V.�(!�l��������0s|3�K�q˲�*�j���q�B�K�7���C3�~Z<P'3��'�|���Q>K��+UԼ�R�M�J�5���{��!��I���&]���>��{r}���"�����L��&�����loe�
� 5g����s(R�~���ĭ#����1W�	;���5����
�۶�*
Z����-3 PvX/��::�w	�����Ų)������߲�yU��|ښO'��va��bm�=��B����j��G=���Cń�߱en�;7G�Ir=�aB5��Nتz�d�]gXN��	�vd�����}h��éMyVi�n����袛��7��ҕ��K��5'-4q�!�
b������� � uoO�4�"p�{����#�5!w_����	Y^���� q�k�{^%{��4�D*]����vcPXA��}��m��%��S�;�Iz��t�&Nn�Z��^�g�x�R������Å<7v-�u�?�aB��Hڎ��*�F[u�1��^D;P�G-���/d,vz��r�&;5=���C7�Hrb<!TL��M�������ν*ѡ��0��T�̺y�|D�ލF�
���������/��C�[��dT�y�[��d������(J��Bq�a�r�VʾE�?(��Ю���nJ�O���#�E�dz"����RvC6���=��)���̛�L�FH~�To��S&V��wܻ�o�4-�^n�N���bnI_fAq�x�|LH��?8H���=ҳBj��>��فgMj�3�'�Eܱ�'���'�׫��F~�x���|6P��q��E���H-;�R8�-���䄂�c�31�"��T��,�3�ᕢ	u�t��Q�!�k$/ �'zJ�fiY_�eM�����B
�&�IOԷ5� �Tx�7ܣ� 8����C�h�,�+/G�R�)��C���a?-F���(] )�W�0Ϯ�O�F~����c�hv}����'O�a1%쵋Ǩ����M������"p�%��^j0���MI��ES5�w͠��/?���Wp:�6������Pr�݂\{*XV�N���%�Q~�I0+�<z�D��x*��&��K���`;j�q1�2Fe�g��\��-���ȉ��_�@��,]A���� �����E[�p+ޮ�A�q�*/A�	3�9K���~������k���?�{t��0��4�״c�d�:�<_�^1�F貧�5��ս#]�Wt^/]�:�j��:��&�%�c��Է����p���|�J��=YNj髄E
>S�}#@��-]2���t�1j!Z��ZY�%@5�����P�O��`��ç����?Ȇ�xh;{.p��mMw1۩v���v8ծ������[�9��@�J����Ǖ!�I��å�&�p���R��LV.\���C����#��\�'�n���d95\��M�����I�h��ˤ$=����=�����C�s �,�G���`sC��q��1�y�K煉�؆���@�̊���	��������S��D���GYh�娐��͏	bi��6ahrM�
�6;�,E���.�$_�ɔ�>9�O*1���$'�����ᬷ�>{��;8��x���>
� �q�=�nFl�nT�t-gK�PQ�l�.e���=����Y:�[̩R�Bԡ�<柒8^���K+}�՛������(Q�F�='�a]�����B�0��4W��o\q�g��㕝[J��(i� `۵<�7��~�*��N�,��KG�����nqۦog���H���?�a��r�uN����1v�*k����B����ë�WL��c�w�_#�X�B����_���ʴ���t$Sr�uja�Q����z�*+{g�?�M��lV�T�W����U^Q��`�;b���T!�O񷡕 Q�m�L^v}ڥ-������6����&][d)�{x��>[�*��yeT���"��YqaKF��%�H����@��������^Y��yޚa�&�b����֑��N	SZm�D�F�w�t �H�]�=�i�W�wp�h���#��!C�U��-q:���#�a"�5$��D{/�d=���!�r����%nP��ܠ�iV��Q��,�T�U���A#}x���݅��Z�Ze���]M�DVb�.�s�i��x�a?X��^��@>w�ew1��y~6��R��͘��|О��+`p��Wη��b �/6��/���T���bbp�
��~�y�O���$5�=5���y$�d�n�/m�B�K�C�WL��жw<E��O�k�Nsg����5�^^6Hg�ܙ�헎W��O��T�1D�O���}�>�֝޶�2y�l�|g�S;���E�^�\�(����������CTի�_��XN��J!�]2�����v�h���]iC�.�Ȉ=����8�<�F�~.�q���:a$�s(*����i��d��I{ݹKHS��������Ľ�B���n� 3������3��T����=;�3�PKfٮb���L��gN�*V��r��]y\Ԉ/�$�-���iu�C�g��+�qٟm)�4��ځΔ[�I��*x�KkKE4�CM��}�Y�����MP.������뗓h���s%����z�8*��}S��zGq����&�e��E
�����Z6`_8�~�BX�{Y[;������:W�yp��Y>������lj6H+ni��	�����T��d̚����kH/A���*�l����*;A�B�(e��O�p2}sy���"���)�>�o'V@
6۔��8�-�ic�%�<E���gVQa���ܑ�v�{$��NDY٥=򿴈O������_�4-��T�Y�V�(8u�܀f/FVu}���a�4lgt
4���_͕�6���4�n�$ro���K�3�ü��o޶���Q�*�pJX#t�X� ��=3S�>[B&f�Z�����EqG���+*Xޱ�6�z��>���\h������Yu�|9j���o���sc�|_���:p0�4���JIQ-B6�AQ�>1�,~Mh؇�c��?���,h����?*	�3�	�/��s�s=V%�i�D}}|]2O%i$,!��>��]�#��w�z��f���)��XRh����t�=�����N�)�nB�u���`B���q�$6���C��;��n0m�V�UJ�:c����@�,��� �Mi4�َDU�2m_�4�̷+*൚��.�?|�7�����-�sj{�lDc��-���7J��7�^���x�2Y4,�5���)���D��zWS��]��ʉ�`�k[tW5uo�����}��e����M�k��QQ���Hz���4k<Y�y���DYS����S���8��E�}�K���S���316��H�P�̼�q$o��_�Wv༞w~$^�G��=E��X��e=Z�����ǲЂ�?�6#C�<��݌C��N�_��q�Yh�p5�i�Iϲ�J�Ἄ&@����L�%��u����Z>��)G��vN�� hA��hL8$��c��HH\���	�\+�%v��4u��D�c_��]�>M�k�B��62�Ω����OJ�e֟�o�'��ZXJD��H7�L��8Re�[�^��ptr��W���gY��AKu��V�����-�X���H_��g
l�7-Ay ��3�u�7j��?!�y��n��v�k��,�Z+�jA�&r�40o��������}�a�,��4�щ�W��,,Ltd��P}���֒�m���1U�O���MJT�vY6Ƹ�9�Of���@�u��eQ��q��V�LYWp������of��)fm�{����[���������#4��Y:FX�ڪ�D��d�2�"�����Y��5E��w��x������U2'W9��?��blϒ4R(<=�s��	���[�Oޥ0ޥ�9n"��/����D9�P�}��������5�Ym�.����Y[�%�)������O3������5j�k�tx�z���^�i��}�A���{%mcz����
Ǯ�_wTXI�f�����-1��5�"�V�La]jS?,���Z�t6	��o��ҝ������(��^(,���8�K�ټ���[�_a}�"f��ǟȾ c�_n� \9$�|���,]>�xݚ��,��ӄ�T��\R�\NT�WL&=A3J]��f#��N̞���xV�LE���^��:�KWs����m��������#�W���F�G�0}��Dp�ppQ�h�;ènf��)�1�Ly�`p�]%#o��U(��E�����Jc���'�;<Y��1#-�O)?��_*�t�{W�2yPK�7LpY)����z�z����W�u��0)�p ���o�}�1�U͋�J�r%t���"�'A�-�v�B���]H�9�{�<�XT���Fd����t��H���m���.^vtGa*�'��� ���Te�q�wC��Y�C�d�&@����7�v�o�.�,��C���P��uv=H܇��U;~9���&��LV \zmbp���w����,��4�=�a�C�t��"�,#��e�kH�5�\t���f�ϗ���.�:���p����DgǺj?.���0 ��ѡe"�o�"�����K4X2��hэtLM���j���n����e�������6`��_LZA��Ḿ�{#�	l͢�y�q��i������Uj�r?F�|�j_�*��uz��y�R�,��b�on����^*�P�+�1�av�������P��:'�va[j=�2��er��!�4�w�Y�p줽�����L�k����wL��n½��ftzӰa�z�4sg�4��A�y�W+(��d�c����︤c#����L*�CD��pFEŉ7��g�.��f�'EQ�����Z�y�Vղ�AO�*�����m5f��B�z�a"����!ޱk*qZ�M8��)����^�����h�E��ꐿ�K�O������A�����cTI<���Ue6��n�ԫ�qHf��n��?9���������hW�6���s/�O4lE9th����پ� ���w��jE	j��E�O��_�A���Z���#$82��	Q-�������&��1级����Mv�����棟/g�̎�eQQa愾����� � ����K����Zg����{ǫZ��5_	Ha��XB�-*�Q9$�J�W�J�B��&�Q(��u^y" �1l����������MXş�5�&��i�8L��LeB,D+�L�*8��nl��kV�씧7liV��/|8ED�q�)������;�14x�5��4f��{�
-�� xW9e'|�Lh^��)�Wg�n�'�����
>e�ʎ�C�amd8�ѭ�����Z��R����o�zT\Q�ӿ��zBoC)g�r>%�,3sy4��%��D-�U`݀Gq��p�A��y���Sh0�`�rE����O?U�r�ax��Y�?��EJd��-�~�X�
kF�/�h���xT3Bʻ~{-�α��m��b���"����m�� ����FP	P6{�!|��ƣ��w��`�ϺK���V�^�b���J���� �.-��z_l��%h�8Ǭh���!WfO�ǂ�]I�w��'�n��Z���.���3�XL�*4�J3ޱ����(�=��"�'O������oWmT��Ce����os�
��j��)�R��K��ϥ�z�am�x�c��>��5����/�K�h1�LM��]~��%ʛi�9{;�{�ޗ<���r}ݯ���<X��1���({]@��=�1�T�B�:�1K�������5q�q�npS�j]�>����u�Y�ߨ���l��L��_�;q�n�8fo�+���ܐ��y6�[�f�*M��yp�n�c���^�x1U����������:U�>r=��w�e>��8&���,IgMm�,m�HOG��|��V��"��9��]������|����
�t�xcO��tR�R�v�����#�J��`O��p�ʢ�%�澡1�&��	��=��+���q�RE?w�b��{�ą���>9��-^7:�>Jy7�},ݠ�|;pD������k]��A=a�i�Oʾ��(IM���i� Ş0ʃ6K�%��_ajm��> `%���?��_��.������XL�[����$�?%��16�>�I������ �.�;�d���,xc	7�F��:m!�{��Y�p�m��%���Y�Qط>���V
�%���`�Å��˃��1��Q?!�p���soUa	8�"����y�]�Ӗ&���sp)�jz�[�^���Ƅ�i��� �OY[��������F��轷�[� D�]�Atѻ�0���ѻ0D����2��QF���~~�{<_^G|Ȍ�s]���Z{�}��2��x�����Lg/F�0�2��7�8�!#Ι�OZTp��0�P�km�arB�0�lb�{�ZX��tr�ZP\[�
����I�v�	нpȼ�����l�B{ ��X�p4F_����5`)i��aBv�p��鯩�N�9��m.&R��2x���p9��s���T]%E��\�4����Q.����K;z�*E�G& ���Mch���W�6뙑�E�*oj�^��˄�Y)��g�i��P��d	?�1yT�00�F(���X�_f5x�]���:L�s�$e*���� �5��ۼ�E���G������HW�C��Ⱥ����u�2�uƟ�`$�T�C/|g}�C`I�:/����T��7N�!��5}'1��XPE���#��y���3�������y����E:����ܹ�"@x{<�z��&u5E��H.�?����Y���gsވйЂ����0��upJ�QmG�y���j!�� 3a�A������6�CڗF���M[�`�F��C���-�
དྷ���
� G�5K��uƦ+����jT�1�\)e�6Q҄���|X����c�i��e��ʛ�H^StE<	i͡��v��DB�҂c6[ I�F9��`v8���U>sEx��M#&��u�@skAaP-��k�B@�����|�ӷk�k5}�n|��6hr�-_�ЉpۖQ.��2�/��-1|{��m��#��];��P��T�R��o��hCܑT�N�-��i��������eϐ���q-���d;U�L��o=+��E jH"�����9�0#II���B����U�����.7A��e�}W$Gx��7g�/�@������x���,���54
(�;L^��!����23���muVyS�ȵ����XA���|�@n���&���� zN�`�N�����P¦R(���x�,�;�8#��M��q�️>˥Q���+0���4o�b��֬�o���	�K���_�=�ц�V�_��%�z��B�t@&�[���c|?���z�r/�������[O�R���R����u�m���{ȑ��N ̮��0q����d��to:F�⃜6�|���6m�һ�<�%6�;��>9wO�w?�-�`\�se	s�/�F@ퟴ�)v�zK�H�V�XfClʉ�˨HZ���C�@(�>�8z��(��yJ3�x�E���N�/��׭R!>ӯ�<a��,�Bҿ�"n1�����G�{��Z�F�s�6�޴�pwK'>/f���m�KZ�TXfzw�8g��>ޘ�q�W���¦���<��Z��"Y=���hB����>bcB)0�9��ꆴ�W���YyO���lR�9�X��X�tY��b��<w@��ʤ�'�ü��m�R�P׶f�~ضv�6�e�w��l`�Vo�w^-��9m=^+�{x@���uv����("bA�w*3U�e��~%+/�2��g}�O���L��۾��S+r��%t*��
X��Q�CT�`��t��������z���+�����G�@j���cx�k��/���_�=@1��ζ��uL�2��A�ލ�o*!�(��ꦑ�|�p;���%X����1�u�?C�Ǔk��@��F��z�����_yV�}�X���O�<xϫmi>�9K��<M�P9�)�(gZ ڔ.I^��b�^,�z����|�eߌ���*�1IN��E�ZT	�0�J����Pp���T�ƹez��6�v��ͳ���g�������/�zl̏N�ἵ��񥢽��~����]�$� ����H����N�|�g�w V�����#��8��?�L�z�j?��0�"�k$B���ρ��]Շ^5��fy��??'�W���_(�!��H���j}����Oo��DG����ʑ��e�����$$�|%'����i��?��L������?�@_00����l񎗜��~ҜNF�Mڌ��T���c��M�顰�|��K���Wh�J}�����M���ٕ�����L�U_:*�pL�s1?Ba�j\l:�v=����!`\�5�₇���>�;�H�-�zTL�����s���¦���8��_������&`�Ě�Ae�{m���=!&��2�ءc�*>�x�wd=Ҝ��aE��u��A��yt�h����O�Q?U2�����g1�(���ȥ0�T2Sˉs�:ɖj�<ۗ���?W�,����s�я�c3�N"r��*|�A��� ߪ�w�3�v�H�G�׃e�#��NW^�!���Z���UJr���9%Q�_7�����r;KeGv,���<�
ie��$�uUej8���<������H,gN-kzX~ze�d��XGcc�	���D���y�����]Yg�3��l��6K&��z+12���t�s�Q��]E�������d\�J"�<��3}i�Ba'�H��nO}��lr�Q&L����3��C��%���+��z�q����}�V"�r^0��AŖ'����^�tw���HO#Oj�SV�O��4J�����u��~dT}�8T��/�`����ހƗ��b�c߼��ߓ��aVBMg�?[�Ѷh@om�lf�on���N���ή�7࿁���^^�4�¤�7��C�t6�$��P8r�����W���:����6]f�v���B�ư�ﶊFg�ow���0'�ϟ��J������{���)�������H�_��r������Ñ��֬�S4k�ҭ+�j��#����t)��R�W��HN�����o�n,*����E�'��MF�D���3��YT�����_=p�z��Ot�E��ȟ��u�$�d��l�)��>N2�q�f��@ɻ�(��[
� �K�&Q�.h�n,�*��u��X8��������[���"�_!5���������+\M]�1Ri���M����h�2KDC3�	�R*+2�(23�!c���a������3�>�ݔ�Do4Qd��>2��-/"��Y��	f8nF
�t�K�8�,;O�ݘT�b�I�$�̜�*��8�O^b됿qB�4���.:?x�\"V"�����!� Hq��[��� �f0K��q���𔘢ቻ����i�L<9�P��]:f�ƃ9"#��%>�{���H�臡�I��1������\}J���(�P�^Ws���dR3'q������dԏn9�<�E(���_��5yx�U�"�OG�;���LW[bF�#�|��̜+qR	�Z���dgR�J�(�o�h���ng�� Y��D8�fF���`�%�Y�Ƙ*8C%�~�@��|.�1�r�洯�]d]��=7����z	��D"���&������8�W��c��щ�1���ǵ������IXi�!�;1:�ϙ�d��Xо�<��DH��VJ�s��5<�N}vo�c��~��Q�A�n�F"ao���2Z�� {GPH@�tp�X��/3�J�!$� ~P�L�����.a��}�o;S\�J������]Oۋ���i���?���qoeD{b����g�����{ݭo�:2_Ry�>Êx)���y��h��d���4?���?�u�?�K�8��L��|A��#4�EF	��vz��PbN5�w4xS�~�3Ҩ+X�~;������J�������#� �
y�p��.L�Խ�)�����3�00��F@I�v���fc=g��}�J�gH����jֱ�kW՘������,|m[��Z��ML��[
� �<m!�u��+:g�-@I�U�g/�*/�������?IT�S[9@��Lg3&FH��G�����8�����o�C�1�F'�I��w�'�h�o�BrG_��pյ��P�gǙ�R�:%�7��$Q�.��G?���g��^����~��{a���'�����(��u��r�����E[4w[���b�W����j�*�	��� �u!���k��[o���0]��aU|1����v�ґzI���/����k�|�^E�Ծ�ˎ��6��&����!�߿�	�;����Q�!��~�L$f/��*��C���(�xD��M���[�-��ǆ�}��JG&��w�ka�*�'୸�o�����~�$�Ļ�҈�@������1��, ~���ڽt�~�&�z��]�'?+~���Ԉ��F�O9��9����$ʙ
ۿ���3̾�*�5}�*M�8��n��r>�Ye{_q���JXc�<��OK��d"���"������VE��6=���K��Q�1,�{����TsA'_X�Q�)ؕ��ّ>��[#��
��Q���F'-�������d�v�B��n�|f�X������Ǜ����Lz�1�酧1����~Pp���e���2j���k�Sl����)��c�h�G�b-y#��G���Gn|�c.(u\��k_���(^����-�[�Oi A	�D76��!8�'�6sHg��̋S���)"D>�
?���#�S:7��e��h"�*yJ/z�2
2{r}���Vv���ЎW��%KG^�20�]�h<�rJ.��>��l��G���j��%ʬ.����������|�������0+ѭq��TG4��:RmFL	�֨#أS�N�;��w�/O��)
X�n�W�+��硿��{K�-w�ڣ'��9��S�✤2��P�PCѯ���̿5SdÞ�
��:�2�_�O��b̍p�ۉ���<Sn���W��e��0&y,,A��e]`_!�{'��f񒬃���'4��Ք�'o�(�l�x@(��sV�g�yN
�O�����̭0�~�N����
Cw�ʒJ�$�LȉS��	��7�$�L#��ܮcc��Ь����p���:�*K����(Hv=^�.*���'�e,w��^�!jX�&�%hԽ���������T��Q������B�[��"��g��1s��V�wB�?z���Лx�U��Eo,�8�$����>���-P�S��iV�.�X�0��V"<�^���7H 2U���kW>��`�_� ��,y��a?��V�p���?~h:�?DY�<�{�liӱ��{�E�����A�(�.X�+��o��竓^B9�iD�	pC6��o���NY���{E}?��\2*�6D��q`�:I�5ì|\76ę)�xƃ��޲�AxNU���mG(�`�p�a�H���#S��-�ؘ��>�|	ǒ��K�^q�$5�-����Ǒ���%U���O�6`D��j�i�_),�~	��7ۓ%�v��(��2����>p�S,���m�s磊C�z�ʸx�R���t���E��,b�V`�pi{��`lZgR�w���)f��I��rZ�H��������n��yTD���rxh-�y�yf����ȇ�� ��A;ga�?���R�cP��e��� y���s��F�������S�(C��pmt�[�#��Ю���N��ʤ��i_��P^�F����>���Ɩ�(�T��I3�~�#����%>fS]ya��,V�ʓ*\����ZP|�ˋAwX�I�"(,!��=�/a}n�Q:X��ܥ��� ��8���^O�|�(�F��y'g��x5�����v�ˡ�!;>ܲ:L����C0����`�.�TZo�"�D:oi��{؀.���a��b��Pzr�8��h~��n��@0�
�Θ���B;��piT*$�;2�|�-:���(SXp�S� �������V`�-�@��;���
E9gD���N�.��l="Qi���m�{�v�>��{�(Nf���uy�g�ĮV�m8��;F�v�I�?\ԯ����qI���bR nY�`������T7���'L�W���%�Q�ӔC�,w��,���y�f�
�F}i�n5��4��(B����QyUd�z^�/WP`����=�T��؊�P;|Bv[�%{h�)�9�k�s0{5�|Tt�4���Y�5���B���j��P���ę~�5��X8�1�oz:r�Pfg�~/&O�63�Ǆ�wxqne�%�,S׻(����������W K��=`uY[]~&��w�2vՓo}�m5\MP�ۈ���|
��Z�h� ���CxG��9ɯ���,_>����a��񬆦�f����n�I���e���̯-:�nw��h�k\��k��&�\����?DQ�&Y_!Ww\�`t�W�	���lA�����k�n��B)tG��\��(�V���z���'��G�l��ןP*t�S�2�得5�%���gگm�ߴ������d���
�Z�������ޔ� ��u�1�������]II�V�'-���A�,���%���$�Om���Ջ��59vNupzE�"Ċ�{�i��F{3�Éׯ"�4M�:�0|�[���0�5�b�>ջ[f��,6D���̜������ ,�{3�����k=�W���?�����Z�I96��ˈ��俍\�Ha\�O!�S�-���x�Rh���I��3�r��egN6ɓ��/���2�摤_tj-}Ox�LBa�'����^��C�p-�RI��X�O����CB�1a���3g�+����E����SO�CL祢��4�����c���oŧ��3�)1h�:���n�N����[������{�Q-Kqmd#����Χ��^�u���[���=R����s��'!���g���
�a�o(vn���[�������s4Qډ�/L���ArU�c]�nz�sw�=�zcyW��{Z:����w�Pʯ^K
.����Z��&��J������۸�1����q��}({�EL�@�[��L!t���t�P��iB��wkxQ��3���KG�SO�SCeL���䏾Ԉ�FgG!�)���z7hRK׋%�!V�6�"�/���B�L+�1c?~͗Q*q�7�#(|�#����` {�x'6�mØ����j�t�.�+�^��?:l"�٥��12�z�:���Oc?;�1�9�u�%&�#Az��{y'���B�����$ ��'�|�^����	������ъ�y�F�kbe�9E��x�{H��C����{�P[-`��da�ۅ�ź^r��p�`?���T�W�o��^�f�nB�-Q�m��\s�4��b-j�mA��!9���n���E��@�[�^u�.F,�ϛ��Y��<��J56ݥ3���_�x�0� �
�9��3+P>�
����{��l�t��1n\��[��a乯��I���z[��26�͵���"�1�r������gf𳤎V���z� V��Q,H��
�Pñ��vA��X�)t��`^E�fy�z����<�<�DT<�n�7���v���$�~Ȝ���1n\�Z�����[�;�c�o�_���t�Ζ��]��6�0Ɋ�(�����P=��w.��\������"=Mk ��N枍}�'�䃕���;]�S
rI���g��wP�g��!�ꃵ�Pڷ��4z�!�S�6x��u���M`)�~L�V¢浸�eUC���w�ݛ���Ti��tN��rv���%�%Ny")ak{R���{U�=�BZ�;�6(�R�T>�u�Y�X�/?)v�{��$ij��هg���kPuK�X�鉴�L��GE���+��F~E�����l���֑�Ͳ�:�� :�Nq��o�����=-|Z˥�,�%Qr�M���8���Q�K_��iEۢEv4A��S����u|�/��Od{�a���7�c�=C��'��vN܇��Ӎ�o���1hX�_��G��Kj"�*�w���
�M����9�R%��s�*�L [xؓ1{�S q8��\�ܨ�K����V���y@|�A{`�<r@rL�>A��L�Pp�����j���7h���B��8n�R���]Ƞ#@i1�sa��۽VS@Ѭ����c��h��"]�^P�y�Pڗ��J(uc)�z$�`�$�s&��`�-qܕ�ʍ��%n��J�/��L�9'����]UT��N!�����xx�:L�:��Y�PUd������Eh��/B#��~|;
�ڬ_���;��`�EM/��vK݆ɲ6�|aP�0�|���@Djf��Ήg�MiK��Dހ�B�E�/�x
FP�[
|�?o%�k����啄��wpC������瞾EM�Ė����;��zZ����+/����}�n=���⫤z6׽�lq݉��j6<�	���`��7d�q���t��J���7��h��D�C3��:+������f&ЪA�x��� �O�g��4C�^�$�i���ti����@ ��&,�]��sl��s ��u�M2���9�-��A���>�2�����$�l����M[��VG��Mp�w�,�Ađ��jI�Z�p�8Bߞặ^>�$횁-�k]�C,?���l��L��1Z�ᳲ�*g1?�j��)�I�m��;��h�T�)q���X{�w�����k���x�!\.~E�.q�.���t$:n@A�����R��O��4��T��m�\#JGm&�p�YT���]��x6�����zM���H
�ҳ+l�5��^�G�g�p)�?;�d����k&�&p҇�DyBḀ#��
fc�;/�ϱ�$�:�ujJ|�N]E6� kiB�p6��(M>���];u �@ --xZ��1~����o��������iV>��i
oC������@'�luF�gj��Q�*��Qn!�V󾐿����IR�j���El�NM��Ҭڡ����HŸ�D����J�
�Es G�y�!�B�L��šy���5���6�r�co����3i98a�/MK����r��e���*��{��u�Eg_�5���t��=����1��$S���
YWjߗ<�f]�c>�AK�H�Pl�~e9?�ڊr������A�Q���;Ρ���]��Q>�	��y��MG<;�еg`�.�������,o|���t�	����-D�@Yaa�;ׅg�<��E/�"��2�*��*J�c��o��z�w*g�2�@�Z�M3������-�2�@�V��Zwh�C4�q�|:0����`����~�{J�%6㏲*2�N	�'�a����f]�
J���SS�v�W	��p�H%�K�׃!�,ND�µ��!9Q��]Jc+�]���)�<����/��Z�
��@{o"cc6�( OE'27�,��ʆ�����蓬e�uN�'	tTB��C�� nw��<C�<�����oC1�{*y��d$e+K���6��W{8��qB��ް~k�'M�A 1�����.��z��B�u7>�Ιs�$8�/߶(�S~��Q���Gs��X=�߆����#�a���L��,��5=O�wB���f���aA���E�tuh�9�&�G׊σ8[y`,��\��r�|�{�_ ߽�\	b��X/���{G��κ�}%��C�a��.g�J��Et/�\�S1�Ѡ?�	I�w��z���R��miG�0Ou��k���֪Q33���}8V�W���#s�V��K�>�ّF'�xlj{'$���.&7���Y'\�����?���o�Y�c�O-1����4�0�(fe�
k'z�	�k���%�|fmUl�����4QP��üJ9��έ�0p��*��}�4"?�=�k�	'��7��P�l�/y�4���$F�ģ3���kH<#@��w�ۖu�Iq"�����I�����S�W�$�H��X�� ��>u��r�,���OF���.��-��7�PE��3Υj��s�٢���@8@h򲳁�T���w��)�KmQ��t���/?@(^�X�Q�;˚��[r�]�z��Y2�"������T����~\��?����D�S	6������	!�KK@��`���j��!��Gi��){�<ƒ�jX�M�.>(���qof+�z�Z����������f+��	��X�Z[?n̴�m�"�����Y:b9�{���v]|�a$��p�:�N�oDì_��.��Ǎ�/X����'�Z����<���OU���� ?�1�'e����(�N�t��C!��g�  �.7ؘ�!�� 1��l%����vk��=�C��5`�pBh�����*Ʒc� �/i����foS�����.����kN�m�~��PQ� �8-@��F-���z��Տ��V�r���e?��վ�&�yHb�u���q�~�X��E�Q�>���	���� k�N�sr�i��^d�g�,����0Q̖����Ex�X�دg
R�f�`p���?��ma"A������J�����yM��Y�f�/>G(V V���}Γ�_5ȁlob�u�"H�@�j%\ۓ8���T◷}:;�bB�L/��e� Dю;]��o�b��R3:T:0������^�H��L����c"h�Ճ��A����*��V<���QJ��ن��'1���� ���Q$dm�]�F��5}������盀��/�S<�C���F���9�lq�#1�_/�����s�e�K��{R�"}���ac���k�;�����p�j>�������UDo�귌���Ǟ�С��4ֳ������ ��%��UB�$�^���Iھ�x:
��C[;�TPŲ�<lw�k�;)�ա�x��)�o���1�{ӝ(UP�k�@U���_z�7�E�
b�U�V���i����O���+a�/0,�Q�������i���a�������}�q9�5v�V@�����$��_Ld�4�5�MU�J��\gl�EKgL%Vg��>��"VY�ʰ=��̦=���w�|��5V��{��T���z#O����8S�L��Lcr
��)�B[��K���5��W ?	�^�<�NF��2ѡ��c�������\�L0�?���a�;F��:k�70<	H2.����a�,#����S@�M�G/JʺK��1���o�S/<ʛ���"��S!������U�\j���TR[����Z1�S���P�W6�8?2N�ÄH��eΥW�t�Lkh$�w�Gҷ�V�+Y�Q�%iò�zM��3K ϿYr�K�*�}y؟����T��uc�qH�>l4z�� ~Sq�hI��ş��y�}~�����a���L��XL�<�U��%$E�l�����g@z'���z�G]RS�JRI5��$ꭗ��$�:>��~�Y����K�_�}�b4v7�M��a�;6Ҋ[9xt� k7O�����&�%}ѓL�l`����)�xKn�hߘ���!m����r�Z"�-�/܃Lt΢����J�����otڃ���hȡ�ъ�T���P��[X���>ha�i����F�B�'�Y��Q:�FL$�����42"��ȵ[�������V {ZL�}�@���g�*i9�4;'��p�m�|T���y�pյ:���m����0�l@R�Cs�ȹnC�<cu�ِӺ{ ��M���b��.�&ݾY�X���h3��^�k�IQ�1$h�F��ˑ*ȳ쐢Ds�׳1%��`�����h�c��'�a/��4�b?R�ʋt�F?��������4��Ǟ�K�q���E�fv��h�|~�0uY����V�Wb�#�A��b�����ę�,��~uB߶�/�;^>�悸���y�8�9&��Q��ɗR��7��DpnG��Y���]ת]�r�.*�)��9t�n�-�vJ0�{nbl��}#DNW ��x`��a��'��]�Y��D���q�f�����!�n��]�Y14��a��Z36�;�6[wfS���������e�#���.��>�*�up��qڬˉ��z=m��y3|%�C4B��R�}D�O�T��	�m�s9܌��>��"����ǒ��8��l���yy	y�����I��%�μI�?I�PG*^_�Ӄ��B����q��+@Q��@��V��OG�/�/����]\�W���HjZ/���&�����,v*��Ҝ.���Ǫ���b-'^@��Z���Xw�8�YS���U6
�a���H/f��ţHN�ޞ3�v��B;�����bk�VZ����1�CS^�"�k����M;��6�HC���Kv���9D0� O�q�Շ��Uè2��V�/�*���x�.����`i���.џqȀ��%��K*{�W}���m������}V��挸x����,"���N
��O�x�i{�#7��n%�BE8CC8c�Δ�����@�ޗ;@��xU![R��:I)m /a�ĭ�O��Tnר�e��k�y�C�y*�N���S���Sc��K�\J��R�w��`��VS%����	d+��>ʮ�8Ȯ\/�J��@�BVVD�&�(��-Q���T������B�"e�����p�:�0������{uAHmP�x�䟚?5F�a �� dW|����H�O������75=�cS�Hqs^�����3.f�͟6�<@��3𞈈����7�ɟ��,�_�Ɠ"�g��Z>�0�[nZ:����������U���u�"�׺�p	5��A�*�j)���ɇ���c�@X�9��}�hFh�vG�0$\	�fq �t���1tչCFR��h���ƲT��m�����C�imQ��5}���j^ř���M?�ڌ�rj2��㈃�:����s��EVH�T7����UUs"_3Da�Gg��mF��9}L�a�7.���]Wn��|L�����x�����iE�@{��,����ݢ�I�|F/�Fbw\���׉̆��_uS�'�1�}���a��I�s�������(X��g�Sn�.���u�y�m|zX��b��/����-�8�ھ�p���!o>�Ӟ{QZM����6��~����'�y�<�𮀝��=:f�G[G��֮��L��Jg�M�&�?UW��񺄾yZI�8����|@�k��ɐ!Em��UD���.���-X督~�����wy!������ޠ��}k��`����MM��!�5~� ��n�� �y`9�� Y %X3rq�K-����h��%��$�W��0�o%80�܎MGTų~�z;2-&�}���G\\gQ2w͟wE\��2i�`+9�2r�w���@k�{��
���>��`�!$����J@Z��c;#_��%D��`�13'�����3E��Vȯ0�K5���i��r{m��M̂c��c�#1�9T�>�V@Yּ`����I�(�7�u:�A7����i%֤���؏nd���#��m9����ى�La�S
c��ZJU�&A�4 �ePy�{���$��<J���__x"���ߢ�r�"5v�܏%sF��=b.we�Ӯ��nz�6����ir�n6`�)�7j�Q?�ɱ��A9ׇNfv��i���W'9�ߜ8,�wJ��;���I�e��2$�.�"V|] 	�~B�S�4,�R��Ɨ���S�������y8�7h������jԝ�Ю[�s�F%J!�9�������ݰ1������՛�]Ϝ��|�
K5�p�?.�P����
��~N��<äm�~�����T곶z�YEC�:�jU��UF/��t��ǳ�j5�O^�e��z�-xN�?����4�;�_?8aO�Ft��\�K���+b�g~����ڻG���c��(�Мls���??�S�`O���g%+y�㛹۰|Ct���c�N�I%�<;�����M���`|4;K<�EBl��-Û�Q�k-�I I� vY�yЬN<��l�����&�ee�)�A��f;�G/9���*ص���Cz=ؽk���oZH�͕ȭ(�I�l�KJ���}Mwu�jkK��K��m���Q��|U`�	f	ڇ�<M�{|���eqcO��}~���y$�$&%�������E�	o�/gg������A2b���IK>꠪R��۩qXҲ�`���`资�qs�h�1����=�m����3�'������ۑ�mo;�ڙ�݃V��K<�ȏW���j��(����1?'x�f��?���X������㹆BϯŐ��^P�%��m�P� |���j:��������w��*�H��Ke�ީ��D�Q�GrXt�i�CD��	��h�+�d��T��3�_���{�`bi�
_�9ɖs8�s6��	�u_~�C��Ah������ō�Д�C�7�4����I�4V�+l8y_�$C_��:�G��O�J:yG�K���$�R�&۫�u[��lqڑ�-�p������PǊ��ii
���&=-K�H��٭D*�^��8�c�����w��X_����1��n�ƩE��ixC�����#�V/�IO�L���_+!		�{/PXw�is6�Ÿe���^�Z;%h���۳㚃`����clF#��I��؀�z=�&5Lw�1M� �8�'Ij�o4V'ܒ�mf`8x�,�^��'eY��9un�L�˞�$�'�#m�n>���)ȴ�:i�C�i���#n�,h�l�~���i%��0��ݩ��N��־�I�V��iq5�H^���]���m�����̙����7��J��n_������;��S�����X}�/ђtg�j�鐩��������3�F۬TcB�xǮ�*ix؞8��)Y��ocRV=��T��l�3'��U�Q1�R��Yz����}¾�f��O��v�������v�;׺.����&�`w�F< �ެ��Y¾�?>P���"�hR�s�	B���eo)�K��=�����s�XN�CǱ�!�9�3[��k�>T�7�:�.�'=�4;�A��?�Ƣ�n�gI������Dm����շl	*�����ْ^��z��N��~	uk����k͈;�{�[�e�����0��rD��88�$��m���ׂ!R�6K�9@B8��:�X��"`����P�^D���d"��w֕���B/=7%tO�#7�
�Q���D���2�!&����:ì��Z;{,Lé ���|�֝���Ǐ�mbmm�q�*�a\ �uV1���V_��|�)�D��ύ0�Ԙ<��k��@Z��������e�[�=�z?��ӹ��h�^�S�*-�En��t�����B�ÒMϩ*�i�'�^���-�������O��^o��<��༶��I�,y��\��ϳa�s�y���i�sQ'���gn�W#pH6�?w�W�m�}��}z"�:�ɴ%;u��drN|�t�\�J�ꦘϭ�v��इ=���[�
D��:�r����B�w`x���e��\��}2nD�ڽM���_�ie��.�'�Ko��w>?m�e�^����b��u����h�Z=D޴�`~x�)�c�Ty� z��$97jx�Tak�Lс=�;���	�X\��G[�g6��v�?n7��3^}�Q��BzP��l�	PF}����fm�ؤ�*�*q���R>���}R�r�Q�Q�8�U#K;�+��z��+�\�P����C:モ�_���ڕ��^���x�T"꯾8�c����n\�J�fM���h�b�M�*�k_a�=h�Q�9�*Ф�7q5,����|Ē�K�@8������*�P��.I��/�C<���9p�{�Oi��,�b�m�[]�_��J����!�mo7��,�`rl���� ��V�0�|�俼YJ�L|��Yu���TyZU�n>��wl�="�m�;Z��R$=�y��-��ivX�E��=�pm��@�q\P#'���Ƴ}�a�heJ�ӄ�oeM�o@(57��6O��w�gva��n����}b*����P���C+IT�+y�2.5��G�}L�J-5lab8b~��U���xtGxK`�r��9M���N[#��5'㨟�_�|�tû�}ӄ�����1��j���S�F�W�
�K���v����C�S�O�	����nd�5F��z�މ�Lは.b;$�t�s�ޱ�K�O-��� ��̉�c�ɮ���{�?�ݎc^�ƅ��'d���Q����{��.:�x=����V[zx���irKqhH� 	ARm�xP�6�(��T�u�]8��1قΆ��w�4��}7��`P�VŁ����h]�A�+,��Gr���p��kR���3������&���ҫ�CH�Td��˂�V����͛��o=iG��ݞK�l� ڌ��~_�P��1kHa�hD���w��4��N�	}�&���<T�U�0�{q�4(���w�KԦ&�M|Qh����::ޠ������3��vȻ���g�u��f�6ܞ����������O�r�Q�*�l�Vz����i~�0���/�ѹ�z����T*|�Д����<4����R�n ��^�qU�J|�|�<����|��Pla(�O1$��7��NQt�����I��f�z\��L^Bb�~�2^Rۋ���X~k�E�)杝�/�	�ɧwe@��ı����T��sL!�G��-fH����*r�6�8���Ą{V_q�-�wYh��`��6n��^zH��b��P��![�FX�t����0K;�Ŝd�w�;zs�6�w�ϻ�C�U�Cjv�{s=j����fk���<ˏ� <I�y��{��q�3�e��1�A:DI#��x"��7;>�9����m���ZW�J������j��2��0׈�r�9������H�V`�g��dth=}�;��l&b�l��#���1��V!��څ�TH�'���K�͔e:�q�����7� 2��`��%v���8�Ş]�:hX�W�Q��D|m# �΢�£@�z3.�~�6#�2����*�#�gS�h�����p�"�U36=�޲*�q\l�;9>�B�~6���#�@�|nqx����8~�W�p^I�̷���i�;)��}��A����Ms�h�1= 4�%y��c��lu&��g�������y[%̒�0g���Z\�c�J�/����?X��jV��D)��CB4�ꍓ ���~�Fn!�X�}^��JF���������zrc�R^��N|]���~'���V����m������QKZ�Z.���g"��x��Mr'h�:ˇB�A��{���	��+�1��b,�i�>/��o�\ބc{zJ*~��@[{���������@Q��n��i�ii�CB�!��-!�� ��t�4�uhι���߽�=���;�̞�3�g�9�>y��/�҄Z��(����}�є^:����ю '����N�w8���Uf;�ׅ����Dx��49��t����^�zؔ{��^ת����t~�{:\8Q�q򅋿�?}7�H�q=�O�Z�n�!A����;�RU}p%�d�?m��͟���z���;! �[Օ���u����)r	:`��P����pqʋk�����u�>��h5͵c^l�.�?:nd�pG�ˮ�c�;;��P�$Ҕ::���7y�Y�0��}.Y݌���B�jl�xȆ�* Ak�rIsb��tg��F�B��Dk�(q����wn0=�����ȽX���"&Ӱ��Fx�ZgH������fw���-�Ţ�
f
3d��Zd}�Y�v�ؾ��Á-��S ��21�	���H�c��ƴ�W$�ȃnbN@ς�3~���W�vm�u����\���6ub�3#a��}��
JH�v�Mn�..�zs�c:
|���<�H%A3�i��\T;.�Jf�������3�rж{�K�׎G�������		X�HbeEDjj�\z���
�Pl7��6Q��2�����1��'x����`���G3�3����OXߍ�����P;��ed �͊8��&wi);��,��9��;����+�E���T�8��~="m�Y�	�K���O�X���x��2�pSO�R�R��t�[ib-�[tد|*wA6����`� :.U��H��s���ڑ�rrX��}D�ɲA�� � ̓����[�8Hƅ��Μ�k������q]�:3	%ᾪQ�&n�F7�OɟW�(��m��S��b��2Є��� ��E��R�����l�n����|N-o=bS��nN������a�� ��=�]t�΋~S��=n���_T�\�乑�(�;1s:�<Z~ٖI�[��B�OOlٸ�b�=���x��	n`|4�?R�Qr�m�`Ԁ���v}���&�ݻ�����.F�.�8�p��N��ޘ=��t�ýTFF�O_T�R��r������|u%�%)�D��Ғ�2� �k��R�d_\�Q�
e,E�/I�H!~z���٧�g���j�r����+���O
�ʤA�.hyV I�ϡP��O���2&�1ʳt�W���
t�JC~ �};�B�/�����˯���(\ع|c.��_X��Zz����mO�W�M��KjNl�:�V�(sc�CQ\I���3�v�u��YW$��J>|�OÒ�t$�_���bM����T���y��(s���h���^�ޛ���ak`��Xe�kq |T�ｽ����Ai�n��!M�ǡQ=��K����u��G.Ĥ�E]�/aM�4�p������\}b ɰ�E��ׂ��f�2����^S�8?�B� ������ �Gr߷]�MHP/�p���rEf�B��o�g-�PcL~SE�k��W�LR�`"�cc�[6+��_���BB>�-,�;!����g���m���f�O��葇16��Ma\F�=�vp�'#�����l\��
��3���=����R$���/^��Q�\�����4IL��N����+��/��Dm�O��Dk̮Ǳ�_s�vOL?WW���61�Ʀ��]�#�����5��;F��|�&�ؾ��������n�x[�'��^�8P����p�C�q���෴���?fb]4��V�������p�������Jn�[�dx�>賊�Os��'+aU}hC�R��V��A�(�ٞ�c=>�_�,�R|�'���c=��C���	������X�ev�[t�B���_�i�&��~�^�'l���ev��N�o01�!�����ߕڲ��=��S���� j�$$ZZi9�����|��
���Z���[��p�S[�f�g]���^�.2|l-ҀVL��yk|�����d����؈�_�#���W��_��jn���7\\/ ���_Q
�n�k@�p�\f�"�9�2C�(���yodD���9a�����������:�]E`n�KJJ"0�������GI���Z��|<KOT��t��ת�-�6E�h���͚����K	9��ֳ��k1��/�nh��Xb�N�PQ�_�P���M�X��F:�_E�};�=$�8�����@�
J�
�:�u���1�����j�*ƝJy�������(��pe $��g󠑙�� ed[�U�oryor&��d�2f���B?�Y�.������/�����,���%tK[�֩����*����쏩�E��V�b����		�D���H�"�:���_���o�g�#��w�����sJ��+��}���?�Oi�b�s������>��S������Op��)1�$c���=_�}�M^��-DT�<]���B��CC���-b��q��Q ��T�ŧ�Y���&q��j�+����<�y�5XC��N�@�#T���mUW1��ڪK-�w��3�o4�Z�e,��!��]�U�8�h��u�[{2�Z�k�^e�T��*����S��s�
Ɔ��$�wJ����`D�S����V-��}Q�l x�V�8�dǲΒ��G��Z�}��E�ASJʒ�暫�c;�![ִ0� Q��s����#�o@sK�����B��h�LMI���BaU<�i�n�&8]�`n���ͱ��=�U��J�	��K:kǻ�d�~k-��~���gJB����dT�!<	F����!�<�IPi��e�!��(�9Y��>�1����gV.hƻ/I�dQ��H����g��i�L�RF�_�r� �Q��[ΟBy�1҄R����DH�[[6���]�gq�H�ְn��������VGDR��5��;Ɨ���AJ���d��r���R���S�Y����b�F�5����eNH�-���q���P��N�g��W?a /����� �p�5��h`a~/1D2��YQ���dBbҿ�'T>����:*��� ��E�w�7���������`���P��{���8��i����h�2Y�{�p-Q�>z��d�{���jv�_�ieG��E�Rq���8��m�&w����|�A�_� ��γ�y1O#q�&��<@on.j"^����
�!֒H��m�� .,t�.W���؆}�ĺ��@{8v�U'tQw�+h�\��*h|�n~���uѵl
�"2�DK5��H�#�]]D)r{� yJ�����0�̋������H��Qi��i�сz4�oݺ�cZ	 �\�%���j&��H>VԬ��Go�8����,���}fq"���2��r�M;�a�c���
��\�I˂[�3EG����96����{���z���ޭ�EHB�ƂSȚY]�1�\�fh��8�|��3+�(�wg�.���5H�Z��s����D�wZ �f����.DZH����NI|'��� ��@���([v�����n���y���g�!�RP=���+W̖Uo݁��-�&�ߟ��+];�	�tI����S�L+h�x��@IdKy�ɉ�m�[2��B�^\�ݫ"�ƃ8�dIl@�-%7ǝs�^�+w2�(;���I��I�;r��y��{؂@9��^��S
����;-��n�{䔤�%ڎW�Ԯ@�����C�!s�k^��
HŎ}J&���!2��t��V~}��)��Z������y�ﻦ���*������R1�2�1j������Q,'j�0�06�ψ�CeA4&z��ιX�J��Pw^�P��}��U��Za�eB�L2�P�oyj<�����q
����]�Ǝ�;_���H��QN�H�*���+H�$�8>�u��1~�2mg+pl���u��a�<���w�����{e���>CDF2��X���I����#ހ4�J߭��D�e�Y=�1ͯ��1��UqG�����|r6�]�_�n��<Y<�l�d�ǻ��&�M�bG5[ѾGɫ���D+�8�.v�'�k`6��U��ci-���ޯ�݇ND���*Wˏ&�^V�'����!v���i%����
.�o�&�n�~8|���Z$!4�b�pU��Ew"��z��b�ڤ��Z���
�m����mI�S�hq���� ��7�(�� �HhV�1���c�o�*�7��
'w3i��ݥP%�c��h��nCy�-��]���=řO?�rn��?�.+��F�* Rg]�҈8_"g�z�`:4*>ѷ�W6'�U�%j(�&"���m���sl-���w�F�!L�.Ba,T	#����)	�$/Oe�fK)��2�����OL�ي����`6�f�0�6��ͮJ�U��s�#��Rճ��!����g���ռG����ҟ� ���uaA�� ��D���I�T�q� �fVZd��t @A�%�t��q�qi���ݼ8�\��y�G�X�J�a���c����Χ��h�T�Tg�,��9�/��v^Ʃ�a�\
���E;�ʟZ���օKSL�Vn�X�JJ 8�m �y$��LY{4f�$�c
�o�-�U�k7�j���s�,��ւӴ+�T*�#B������H�@_�N	����{��C��E�^m)Ǒ�Q���-t��$�=��Rz>뗋�N{ϥ�$�ː�[�U��:�;9]"���Ii˅MSiL��X�CT����J6��"0m��=@�	�&��3���"P.c��рQ?��׫(⟷�"�9�låT9�bf�4Z��gּ��ݫ,oG���*��2�s���]��&����^���B�Ē�̆!P�VW���DХ�f<�4�Y�u��n���a}�[zj��s���pdb���q�q
;���
�G.V@bA�sv׍��sR
M�Ii���!�Y�i���˪e� ���[��{Z���W�m��/��U����UX�)�>/�����k�,0qH�l���=�Īq���	����9��O����o-~�{�7��ʋ�{?+�]��{<�!�r9�]%�l�'�E�v�y��p�ި�z���`��3�+t=��tX���F�)x��L�)�@�5�1Q���`IIp^5�g�2�`"G�����C�ǤxZܶu6+�?�Tc�dp�ZWT'[�	vՙ�)7�~r֓<n��8?�~>��}��
4缩�I�Ĭ*,Z�r#@�zX���[K�l�_����6S�|�]��=CE��nfZDv��m��Q�Bu�c��M�r���Tҳ��v���͗C�av��1�N�r+�C�_ۓQ�ڿ�&R���i(��������7,���Fw��ZK�RqR ����4~�G�?���nDn�~�����3�ɨ�hW R����𬏶��o���� O��T�	�<(��!�iH#i��>gJEw�� �)�����,��������l��S_�qԔ�B�l4@�O��*	��r3I�P�l�=�hB��:�:v��jI��~<d��o@�ώ�/9���Lyɶ+B�A�츒�51�P���^�?�<p��;�V+5"�i�C�aa77�jF��{�#��C�����Xq眮�-@20Fz��iO���.N�C�"oǬ� ����#|����(e�h��MT~�K˨<942\;bO�"A=�V�fh9�Qe�ھƁk�*C.^}󂌰�N���I��!q��8�	⌟�Rv4!�i���e�n`��l�7�[�/����"d�!$KczQ�w
��I+���z�E���)������R��Lw��2���'>R8nϛ��>=��Ć�C���g)�ө��&�@]���ќ��������c&&p	0䢙K~�Pg	G/����B�S�JQ�(/�&��X�J���&�9��A�ȣ�4��=�����&)���&�C�1񖶽���2[��ŧ�0f"��!��f�3\B�<e�vH�R��W���wr0�ս�,�k�3���e4À�
�2�o[m���7*�W}ԝ�ӕʺ��l��$��TS6�KCG8���y~誂G������o�N4(���'- jB��*h�B���	���\�#W���yf�������3�b����D�������ז���v�J���&��do���K'yȭܼ�j1���97�ؑŤ��z�{��jU'�/��8�y�$�JK��J�[|\�<�X�o�s�H�-B��~E\eA�o@��m�1uk���-Q����f��t�3�����
�~��{���?=�ί��'���~�y1S�|�ɔ�ǰ��+��K��+�7	��r�Ә��YK:�5v�|�XLiZk�Zi,v�~q�=,�C+�O��W�;���(�����z���]�(�
�sT?U�y�s���:���ID�%�4��ifpF|���|1��BT��`��b��!G�y߷��-T��GrT��N "��,r���3�l|����o�`�F�4��j�%<���0��6��>e���o��M�i�>��$���0Jz0)��,���U{��;ͤ����/��(�g����?g��N~2!�5�T��9ڈX��:�E�4Õ"��m/��zd�o3f�≮R)�0AB{k���ϥ9E��-AyQ��gCOa�?Ia�RI`wF������S���No���Jw������
��o�z�7"Q7M���^x;L^.(�%��������l�,z����ۨg8���\�i�R�׵��&�
�[>z����U[U�������_���]�=X�~:���[L�Y�}�Y0�]a�k��N�X����W�?II�<�zKp�\m[�l���J5������sz0��aC^���ӣr$hg=�!�B�Ͷ9�!�I�q�4�[�0B�I#�����E���Z:���l/,[��|\շ�腑m���x�<x�����p�����s��o��Xh����};`�":�"2- ���Q�o�ק��qݩ���5G�R+tz��������B�_�ӱ�G��H��_q�����e9�WZ@�]�*��nyj����M�.�t�+ypp�%�y�L�34�߮T�luI,٤��<g�����v�,�&��Z����#��w5J(]���\����{ɦ�cn������ƒ	]�=�ʷ���pOI��ZΗ��������?nA���3	\�iP|B� X
�n�:�H"��=��_H0j��Gfx�q�w]���K��\��j̮�1�zn#U�y�sO�7���[�H:4;��/���qՁ�x{٪S�Dp��`1ۙ��կ��&0ӳ��ȶ��L��l٣�V�9{����ն��Z��!L�`���GBF��V��j)����}��D['�ӻ{'��Y15�mj\Ŋ*X���	��yo&�\�g1�����܏f
��>�q�����#|i"��e�Hzn�����C,�cGC����vs5�1�y�����'h�Sci����j1���l�c5W ���Z�)C��j.9V��R���FV	k��H�>%>>~�g�
^�2��I�G�E��7�Xc����g�tՎ�?�+;�������ʲ;)��	�@�F w������pA�Gne�i��h��Đ�Z^���p��v��:���q�yT��2�KV�W��w��V�r7�pt����U�����f<�Ј?��+0��۝��ǃ�7~ O�/���R��l�R�z�;��(�^�$�4R(�_R �ER���k{�Mݴ�MRՐ�B�.)���	�a䧴��!Dg4���n��"�.G�O����x�ޞ�Ot~V�= 0"���g�9�>��ɠ�����O���>.=�t����������bɐ��U��GD��6�a�4��E' �O%��Q�^pu�D(b3����.|fPH��c0��;���\�	P�i� )�g*�%g��x^ȴ��6Jͺ���I��L��?�9S���#�6YL��0* �Nٷ
�<��?=�1v2�HMx��#i���II2Ĝ�� �;�$��_�6���\m|�)w��"�>�`w+w=���n��^2Ͷ�y�J��0׵�!!��lo[@��������P��>�t��^�����h�4�y��_��-�B�Ռ�t�<|��A(�+�'R��EQ�؀�d�_�C�����������䐝�z*���ۋ��������PZ�+	�LlV[��G��ZkT-��i��d�'�#T���r=�>n���N�����H�C?�_-~/ޗ�Y���[^9P'?s�m.�Ly�."�XǺ�!�~��8Hz�b(C�B�?S�	��)0���h��X�ru�!w=�~������,��tP��>?]�p3�*��`e44*��mI�c6�0Y�-�K����$r�Y�y�	�����Fz���,D�:��*�HZ�"��z�#!�z���FjL���&�&0j˳�����~�԰���D���Y�C����m�.[Ǒn�����F�Rm� ������$˓�zcwOQ?���G\ ��E������y��ߦ�L���;A>�qi��s������)d]���j2k�;�+�G]+=6��q�H%Ad�m�E���Up^ѷ��F��\���X*�����"�n��%o��h�ȑ����?|�ՠ:�I��Θ��3u�_�%�K]���m��-��2��<�;067���aბ�vz�o�1�WlrK��f��h��j7�����$Hۀ��n�A�b��(�Klk�m-��R�g緷p�
��u*��"$����Y0$�����gᄜ�7e���h����1��U�c��j�rQM�ޑz:�����9u��vgy�\��|����A��C37f���2�u�E�H�W�4��d׭�3;��&��עl�q��(F�B����?E:$��v��1���Z�ǋ�;�Yҿ����S}x�c���v���;���g�xd�R��`몇��F�E�ѕ�S�*�ɿ\��G��GS�[uz�M�k�d�G��c�kdL7��!>���+�ʨb}�wX3��	�&��Ť����F#I�y=��}'nk��~1���N��v���G��I�Y�kջ�ۈ���{������V�?I펔������V����9���i@�	��ZC⁑�S��7�W=4=�d��+ɕ��+e%p7n��&ۻ�8#g -ᒌ�MoZK��l[*)��Ѹ7
�\�s�)D�K�+�^p<�����F;�5��K�V�k=M���o+���-;���gc�©������+�U��&,!b2F�2��S^�;��Y�?N���Wې������H���3�ދ'�p,/�LK�v�0���x߹?���bj�F8�F,.U��W�#�	�.O�I�6�;X�N��Lo�<2��fVmI�\f���� �'c	3���r��A蘢c��kb��h��c���ah�'��!&EB��O�����Ӣ��$�s>������S7��t�jlTHJ��֤1�}�I1�5�Y���ǚ���{W���<��EGL�mr3W��ͷ~��J��溿��ϋc���m]��-�d
�:Y<���CqP�v�7��yw�#�NZN���EQN�J� �Ba���y������X���o��u�����9�x�&v��p 'H�����7y�X���qx�x�+�U幈���5�v���^�(�$r\�E����_��}�a�Y�ȗ����5׭z�?�)�������~���g��u_���B�RÂS�r?(��T�_�nF$����0�}���$ve��듛�=��;���-�2�P�<���.红�8���3)��r�0�K�=Pm��� ��:��6��|xZ�ď>�+W�V�ȶ�K������9�\�gq��ij��]���^��vc��T�b-�b��i���I"�{����:DZ�x�M ���FjJn��l�ku%̚����mt��1�B�2(:\�T�pż��z�Q��-��p�MxM� ����!^	���ꑛH����1r��QDTf�,����j`�eF�9r��B�\d����PE��.r �ȣ^F*qy���.�(��0t�n����K�V�F��#�w����w.<+��;~d�n$�|�wck���N�y I�m�`v���!�@�^��`�W�VX&|���}mJVԹ��GO���O�jD��ӓ�$��$�4���p��P��d�P[�Y|�'��byRY��Iu3�>��:?�[�}P~�Q�	�K�V_���3 �F���U�Nd�Fu{`9qS+��@�3�S��s��bq~R�ц��k��f����8n6ѯ��d��-Os�kJ�P��ŉ�Q�T�a�O:�>V(��T�������\�jE���i!ΝO�� �_�svg�w���3���r?�U�d��aNǾ��>���2��{n�VᨷEz�~@uRT�n$C����l���c,��i���x!w�J\HХȿ#W���_+j�O��>?g l�!��7�1H�0佒Y�à~���<Ќ%|j �w��e�niG��BKЖ@Q|I!Su�&�¥���MJ�g�
;�F��݊D����P��Dl�|N�����T��q��nd\*@ǂUwj������c���͜���ex�m~6~X�P�^���qĕ�1�[1a���7-���~�f��.U��ǒ��?��K��x����^��yq}dJ,�ܯf������_�����%��':�5�uO���}��2V�T���ВʩC��h{'��↘Ǟ���h(!5��[��[���L
&
���S�0hT�-tرlIE��w�Ļ�8g���r�<��{���Qޗif*>H�j)V����GF�	�%���9*�q��ڭ��^�*��u�`D*	�ԯ �*��J#8作�G��H��*��� �;�h�8ܥ>ɒh$�]A�WE��Q��p���?�cʊ�VZ-�0�N��k�Ô{��#y�:֋�y��=G��s!�&u�/�c��~y�������x��Z�r;vet~T���+����|����F��lȴ��&��,�|�*��訤	R6����`���g�L�\�;�ɟZ�P�;n[ ິ(۟��K&�S������<�m�Nt�T&��AZ75�0�� "<��7��O)����ؑ1�v{n5MvfIӉ9ãK����?G��}�E���  @^w��kd�8��LR�w��zf�N�ٟF̚���Uwc��.Bȟ�uY���� �ُ�BD������J�B�Z'[��A��-�V44�������V�׬~�K����9Wc���'�>�əa���Q�>s�M[���YZ��Hc�B5Y�������]m��V�g�����aڇ�����DP����?%n����吜>鯝Satu����Ԅ?΁#���A3�0����&dn�@��P���أ�M��F5�R��X���p�Ò�q��藪J�Ā2��K�ӭ~?X�g:�l( �޻�U�u#v�o����%a��,T�ʐ�=�J���;������*�E�������;:�"�e*�}�ֽ��}ߪ�%�z22�A��X�(�?bO��]K,�&��$�1�rV��\l��u$�pˁ>o}&V�SQV��yV1N�y'x�^�g&��4)��s�P$e+Ǫ�#@�$,/3�#tOc�l��b��÷���r"��/%�J`֠�E���'���~�����[p*	:�Y��L�h������g��{0fp�0�WC�����*"YU��k�LK�W���l��2�~c�k8j�	B�ڃ�氱J.����^��'b����,����47m�B����D�͒���me;�(��4�]�5:��C����{u}�g
�¤���(4�BN�>�8s�I#��5B��	��:�mf=�d�"X<̵*XU���F��{aK�^`kE�%�-���6����S�{�$�D�O'��Fhqe����U12��f:ٯY�ѳz�*�8��~�Tvx�~��e&�[�%��8۱���EG۫R�O�L!�MV�~��x�� ���u&�?���7Z�-�ߣ>gm�6L�PH��p�R��xT?��3G20��]MOiy��:�h����o��p�r��j��}�p)��fhH�?@&�>*g�����L�u���O�4�ґ*I�r��'қ#w1���
�£�x:�+̂�A%�=�w����{~��E-=w�¬b���C��Ȁ
����Ӳ�	�P$��?#���\ڔm�剜��ړMz�ZN6c���s�n��ӭ��7�tVBXn� Ǵ��{/W���8U���ؕ����s�7S���*�n:4�>0�،3��S�t�Nx��|��	������V�QTx5'�!B��G����`��W���!���������V���p<��F,���B&�DC�C\%)����Qr�W\�7
�n��d�PXV�#�ŵ�Џ�؛��k_��mF���ҙ�
�x���Ȅr�N�a�M�AR�굄��т�:l��R��Q��p��+A�-M�
r�"w"���Gc������ɋ2:�;����.��Iay�x����E�B^������&[��cH5�Wd�~������5���ޛք��5��Dr�����CX���p�+���\$�Ë4˘����7F%�!�iX�4�$��3�)�4�Z�}׆�4�`C����l[o�cq�� ��=��B�`1B�~Ch|��(���US���]���׬����d̮\����z\W㐒��+H$�>n-��������d�s��p��s=��ֳn\v�ᤏ_*I��NI�MX�����(7��F��,�V^1����M����Xv*>����j3����xT��`WJ��:�]�ѥw�O��Vx�"�m4�\|g��x��t��5�/x�_m/��6s{᫳K�8�,�E>@C ː1�4n�w�7���_�%6���u���j2^����9�;�	*����fi(�: ��~���9�B�8�I���6�7��оƂ��w���|zؗ��;P(VbX�x���A$=�d��k�_�Ѳ=����'�(��wl��!L��v�5Z��3�Ԛ���8��K�i�_��{��́�l���!3�H�������R"� e�C� }�(�])��c��r���G�!�ƁL�FҐ���8�9������Q���*]�:�ͺԀC�E�v�E�_��-L�SA#���5!��*��p�{�����Q��b���4�p_e߹N���fq����%S;�d�G\l�8\�B�Gìk����/��*�ѝ��=�0ky:Z�S
d~�ě�S����򦝍��ȑ���T�,q�Y��d&�!|�1m�r��}x�OG[~�[��#����(�Ђb&&�<:�<�x<��Ҽvby�2Q)��U�2F^��8 J.���x+s#�w��Z����>���;�T��ߵ�q��ex̵��	��Yi�(�|�)uD�C!����q6n����2�O�saP�c��ූJl�6P���:<�3�3]�E�rg�l���N���������y=HpO�d�!e�H�i��D?k���ֽ��rY�l��o�N���c��	�gC�m`0)?UAa���l�������f�;����l�g�"@��f. *K�uoRJ"/���� $i\F�����ᾟ���3/1LϺ^U��4v�D3�\�Ñ������A�gۖ�[���wQ��Eƛ[�'�xId����p]���s�R����1��_U�Ee��N�͌�֨���|Mw�B�8M��֢R)4��t��{{�����<^���9�"�������W�a�>�:&i�F�r���4���f���Y��;�ʒS�-�L��r��c+#�u����҉l�gfٜ�O��mS>x��F��7�p��_�Qa��gG�*5����þ��u�379L��ؕ���0�KO��c>���2���9�� �#���ࠪ�jAθ������w~����3�^/�����)�0v �N��r(]y��N@0���U1��vܵv	T�X7��ak�@����Z�Z_����I�!jhg[�c�K���*1�^����^NBB��)�(�4�N�����Nc�Q����.i���Eap�N����2�|;
�]Ɋ���������;����^AQ��̜����E"��L�G�)ʛ>������0�gl0��8y�َ��{����Q`��R�_K�T�
Z�b�E^���<��&u��s)��.p���O��>d*j��npq�Hs���~ƾ�J�LCG��K��@�s"ȷ��ct��A�У�޽Up+=���pīc�������Z0k��#&$��-M4��o����6�uo�0)�6~��)-�{���ů��`FvLr���摑��}4����F��Y�D�8#�~�܂6���U�H���7D㞆΍fM�~Dڻ$
���Tz˫p;�&��	k���U�g������F�ㅡ��Њ�ǓI2�`?l�>M��OC��;�l���?�ˈ��q�����o9�ò�����5��S��no���~w��B��*r�;���a<���g $QZqd�qd���Tb��b)[_jp���&c)��F�y�%Hlp�c�����E�?�Ov[v�zO�~��xbi�ٛ�������#���a�:S3~��Bg,�e]���K����9�) �T�A��J��S�P�Rk���8�6�^<:/�in�UO+�>p<���4��G/��.�T�\��|�R��R~��bTى��v������!���:L��6t����y�~�zMuf彥�=�ؗ�F�
8�����pL�q�R�d�B9el6��ܲx�9d�"�y�7�my�6���cD{�hL��={�8�4Rϼ��ђS��T�9 
r�w��~?����������_��Ͼ>�1�O������0�T}����d�@��0���ͩV���6J�$�6��;����T�f���!VS%�'%I�љ�{q�k7?^����koΤ��5��"���h�p��Djҵz��=~$'*��/�
�W�nf4�����ρ#}�Ťd�
�02;1*6��V���>��	F���5#{.�⢟��R?^z� bs�-y`��S���]^�]�Z�p�s��!h��ay����m+�R�nB�x����h�́�mu+����o���Ue�ɒ��]b�����Ưτ3��]7�n���ׂ�^�B��33��F����r�6WQ+��ȥZsNJ��-�=V�����TT��Ի;t���ߥ4�M�B����K�I����z�	T��O��:�fd�׽��#UHmN�ef'�IU[�>�L2譺��5ڄE1���S�Z��\�C�#�R��i�9_'Z�;�}��yh����Y�#��I9�H�O���pc���Y>�ʆx�.�S���7�5_.�{S��I=�G�=�&9�=o�i�}�J,7s��zR< �����Y��� �%�J���4�됐۵�PqK���������^�$���I��k��+��U@W��_nG�՚:�ۘ����'������pU��o�`�\��$g+�����X[ZO�!6�0B���m{�z��g25��Ej��S�YXjz\��)gE;��{�����q8Z��}=�Z��vږ�a-���2�e��ݯ�6�Rm�m��-r�_]�t�Z�$��Jhm�:��!]���@>���5��Pz�NSe?g�a�J��Z�jk���-�������ԋ!r7鶽Z(޷���m��,�]���n�>2�JtoΉg)K��!��Iӭ��P���Q+��
�W���ޗ��̋R����WoWS7K�Q����Y;��e+�!hW��s��;��ߎ,�P]�O����i�ёym�6����E�xD+	�m�T�9�,���>h<�\�W d�Te��	{u�RGOſ���Vg���J��v�'�=�D���~���j�"��Z[��:�$Ж�����n��=z�遆Jb���[;U�U�/Cc�i���i2w^������ܐK��,����
�dۿks��
G#&@'�bp_5yE*Iww�	��xx���eC��I�T�_o�u�ܿ�8���_�zԇxF��Ξ*��k��k����9�?��0͚��9�c?=��_��=م��^�%f���O�|��whY����XP��o�^Z�)މ%-���w|}^O ��0'�$-��t���v��"{5ekK��t,���5:5�$ԑl�6��]F���ss_D5�-�%�e�uĜh�o��b��d&E��y_���+g	oݬ����x����s��z�/���h��gܭ�	l��r�����8�:��H@�:� 7�5!;��T�eOr�u�)ɉ����	-6� 6�
d��!�'�=�s�"y��t�?��ppG��[|"J'�G���+�����B0�
���M�a_�0�4�~p��(��u���j�q\o��bB��:Ā��H�-�ַ��E?��8f���>w'�~h�{�q~T�\7=?N�^$.�����pI%�t��O��t�մu���$C��Bj�����s4M���C��C�[����5�5��$��\�A�Fw����}SW�>F��������d*�����MS���=�F^��Fe��Ee6�3�N��[��Ԡ�9��0M�M_M�j�?i��'�8ZWX���c􇷿�fϦ�JH\��(���"���w���-R'�����S*|�<a?�1i+��4�l~!7�J��B_,��f��ڞ�,��|�2{�R�)��zk.��e��Cv����%�S>-u%�/ �m��z�3`c���C��!o���m%N�wKAkuF� Ǚ�K�E�����7�?\���D*�A���!��� ���	w'6~��<.n�퉳"'g��Z��B��	��N(i�|�u��˷,�p���|[e�GW�����S�5�_�!��3§u�r����򉈀���堺�r�w�Gi�)���Îw�x�ɕ!����NK��6����׵>��ߜ�,�o}B�En����<Yq:��(���������U���H�u��p�'<j}�c��|��}�X���@���Ӯ��C��q�o�̩TN�Brdi��h��%�D'�ZF�)-&b�
�����6dIc��3���#��x�g�������������1�羯�{_�������~���!�/��?��x�+K�ؿ�mS�~w�ɚk�yw*v���}bbi������}��UtW�;yc�c+��'ϳ���فj\�F�-��N�Y�`3�x�4��l��5G�_�U�p� =w\�q��)�W�.t^U^k��/���ɷ�7>~�}rW��򉥖UF"����[��p��5�E -&��s�]!���T~3�Gq�"���-�C�l�6����FJ�>��ZL�����+s�djDe-��\m0I�`}xJri-m�3�$�#�G!�]Y�{K�˾ֶgY�Ɲ�{�]w�I-3i<��P��<jU��j�v�����������A�Lݵ���C�/6�̘�s�0XX�f����;{�m�F���՛<u#�T�[PM��mn���'|�'׆���G�7����Ǽ<t:#�e��w�rif�^� ղ���ë���{�˕�c�?d�����n��z*�Q[���+�
�R>U�]��q��@�FV�Xg(���(Q6�ʓ@�Nl�2^ۨk���_���j�r��ɡ�^�+:�5&�iJ=�ċ����E��m�z-�����k�C��߿r\�i�w��;@�����U�;?��:�G�T�q�H�a�>;ʿ)g�+�[��g,q��ȹa��͒r��,�]-	pX��(=�;�#h��K'<���3}��_��Jl^$���8TL,a9.���
!'��{�d��f����u���;�*�V��=L�~qP��9����� ��7�}����ܐ]SknҎ�};�Z��ĭwD&V<�֎h.%6S�ݔ�[lO�3��}K����1��÷HOJ2�I��K�0=�-���������/P<(9۝;���{�_O��tU��J�D���<\Ӫ���	+���Ap����`V�y�8? ���~]Y��?)fWn��_��?UlEW�o�_�1���թ��m,���s�����NAٱ��9 	bM���ŌC���hh�
-ߔ���c����ww`�^���B�r5f&� �5h�nꌍ�e� �[�,��N�Z����-?�u4�l�؏7�@���Q������|�wl���n��k^�����������׿�9YP�=�3Rߌ�w�]o��05�7��0Oml����}����I������qIΤ��C����_����;ێ*��'� ������>~�Jm�7m��µt��y�PԮ�3�ZcAc��h,д�7�{M%����X�!M�����.��HlU�M#C��rǇ���`\��Ko����fCq$�3{�3)�����~h5w�S���ؕ�.��M�a`����r�s�p��#���z{IG����v0�̽�<�F��~�;�.��?+s��wsv^���U��{8�l�|�J��c�F�#�W\��������ccbY59����]G�ѼNRU�6~��B���u�dn����Z��olԘ�@E�['vϞx��^��[#P����?��鰰*�n�0�^hc���(��=�5���H�LC��TØљd����T�Iqk*�߷]-ml�m�ƋԀ�)��~�!<��eih�"WUuTwE��<NYH��2-������9��KՈ5�q��e@r|�fKc������@;|!t��˧gjy8�q����t3B�mnx��d������o�Z�ƹ�c��Y���~��k�1�p@�cnj����I�|���a�3�d+���#�էMe`a?:\K:��4�Ȇ��G\�?�2{ 2�If���s�`(�O\�Q�n7�����m���];|�o>n��	?�����a&.vs�ϡXs���ą�5��K`�Df𭏛��������n������
�)�5_���/�,Ɇ�ؠ3�W~�$^7�e͙R���eo�a6ٽ�E~�(''G�g���*�|ѓF� 0��pXhEE��ß7�u���(���W�t<��:���ou�ʯ� ��7��ל��r��5���'���<�nJ��n�<k� ����y���Ʒ����c���t��s�����\*蹗��0m�\��H����x��h��g���jM�v0�%��G��{��`w����7n���G�b�zb����8�A�먪�\Ǿ�Ɗ��˷�\���������I*�K��a�տ������M;Q�~p2#��4�� ��J��o�'8�x�N)�
:q�Ϋ�qi�U�X���83���t:�U��n�7en���� ��eoo�ɶs��T��"�1����������(�ӂ�[U��_���Cl��K�������z��I�_�����2?bzze��2�z��g���'v(�������;�e��Zs���X�����~jz�����*Ȭ+A (���}�|^�H}4�����;*`��AN�U���Ƀ�x����=0�~��_�����G mbbW���bi�]]1�΅�n��Ae{�<y!�9!���K�$��O��@;\�0|Jbb��O�X*�堸x�i~e�A���6��z��e����S&`�<�j�d�u���-�������ll"��|U��;���(+��蜛�x��<㨅̜��Jc�eJ����F̲�t��mۡ��\�5����i�&�1��[ V�a5]��$��0��T	>������Ѧ8��Np~!��א��_��N�0�7�^���А-�o��S��k�i���
��I'���7�7
����5-Fͯ�XW�������TN�,m���?��8�OS�5��p�R�5b=�~߲��}V!�%HJ������`�9x������I��)��2��OV��R�W�kOI����Ѧ�P�����ڟZ����S��^4��4�Q��R�������Q�g��ϔ�P�;�_�'��kO�LƮb�ڔ�u;Η�����f�[k�L�*7����̶A��,��s-��r���5�ŭ�7�F�I�<�Nb6�":^�����h�6L��D̲��p7�^0�^-�H��6_��Xj߮�"�@P��������-�(7�,�2����D6��������->K@���p?��P�w#s�Jwf�ݫ���}�UV�a)�	���oj�kMn�ga����`
��#hdg�Zyy��^"�{��l�\�&���s�)��&���A`�;����3�v�W���ZK���8��͛s����r��55�!�}G�-f��{l
6��|��X ��L)L#�`w��M[C�XDo=�?�mK,4��q�a���g���,�)ا�;�>jYe ��n�#��E<��v��G�̧
xeX}��'�13}��)5���ٯ��现p�/� ��}z�����o���:�a�)S~�:��-��O�GR��˜gM���F�K�����R��|�/���n��|��nН`�׿:4+0<x���b-8�T�:	S�n}��~��P@-�`qO!VZ����1��F{�lq���{�������3ޣ�:��?����C��W��;�]M7C��vk��%�l��|�h�mwU��U���Ƅr�l8ʮ����lP�
%ݖn��)f�8��?����ET}�;�p�Ǉ�������F�C��(���I�&��j�e�ڟ�+�����=���V�#=�%5��	F�g�Nl4�X�o/��z��R���޻#?9LaMNfj�q��r}�/�f��sZ͵τ�f��Y�n�T��x^�<�!�;x�m�أ��ع�+�w����s*��_y}R��ɻ��+{o�u�T�Ӧk�B4���]ޟqܚ��8�~��U]�(λw��]Ӣ���s��٩�Z�O�E?)))ǙE���g6?�Rw��W{�;~V`�2T����|�(R�p��B�J�j߾���=-NӜ�"aH�d*p�&�]�8.�#Y.��ݞ~�'�o�� �Y�h��)����#��ū���זfL�,�Y`�����/nKY�֙S.�am�t������v���4�g����G��~	����d5"-n~h�>�"��B�y�k:��j��!e�/�[��Ԕ���-<wͺ�#wq�{h�=�TF�e8'QA��E�C���k6�1�R�d�am��Fe����|g<���9 '`���8��8��k �J�B��*��)*Q�F��mm5��̓qy3?�2<�K�+�2C-Ε��c��ܩ7J���q�W�Z�s)mɔ��qim	(���h:��c�Xܢ������4�1�8S�4�3 �ǟ$��z6����̆xu��&�4�����.�SQ��6����I��ϰLa�z����$����;ߞ��	�Y0ԑ;�����![86� |���ٹd�왉��V���)�E�Y�i��2��BP^�����w�T ��ѥ��d"�gJp�4�L���OP܅	܌~0���V������u�Eu�wz�ީ����4�
��w�;�@�;��2�Ǐ��������Kzn����P1�	�CF��'�G�}v�\��������5�5u�Τ��V�����C���(Ͽ����i���u��#�R��V�)�Mm���'�(�M���[�] ���X���"h*��C���q,����2�T���U�ԙ��,�^��0X�Q�HG]����n�ߎ��B}�Y�R��J�9�����Ͱ<ȕ�DmҤ|���解��NPR�8�=��ř!��d�����a�֟#�ue�=� &Xxˏ3 � �D�]G�ڋVu��R�l_�����Q)h���x�F�π��s��<P��&觃�;Z
O��L�d�
Wo���mAk�����r4�U�zju6�ґ&�^?��X�� �>�E��$�p�>�DX*kNm@����v��oX���ҷ0Od���Y����S��_v�t����Y��*�Pf�x�\���!�ќ�	Zk�3ag���پ��4����o`I��g�~��~� M�mB�F#��"4`���mr�G�1��J��Us�(����8�<���4���샱	�ӫ���l� �g��)S�Z��4U�j�H���Feҟ�=6-aH_�~���䱏 ��<�`%k~�4�ۅ~�;k
�]�p���+�kw����lh�#�o鎤H�Y3�H��	�H�<uXx�{
Īv������MI��k*o�J֎cB:��i�\���_�<	��*@y)�Q!�E!��5bU9 HR�[�oV��H�:En"�`^[2�D��I3�L(�+L�� /��-,�����	�`��~�ⷷʹ�Z��St� z-�Y\�>����Џ�Կ֎��,=#k�!�0���lb�<@u��p ��$o����H��fĕf�]D����no�ߎ���M�RPA�6��������p�'yb�=�����(?��������^ *�@��{!����D���,W�e���}Q�J�}��n���<�۔��샲j˨~�1�7���Bɉ[��
N�>��<gD/L�'��A�S�3�!�e�D��ݹ�>�>�!�����������f��s	l��BG��Ë�Y��<п�b[8.�O�d�r��2b,^�R�-(�B�I�O��d����4����g3��O���WB:�+��i�~0	�����;�8 ��͸#����l\�싷�J���O�`����CDFʚ��P�qX��ky���
�jUT�� F�'�^gE�l�8.��f#����d���+Q��
gQ=@i�/ތTw(%�
lNN�j�un�iG>25�d{6�if�G�OW5n��N*�%��&�g��	�DZ�@����2��7@�r�����a�Y�2��i8����k�<x6�m�H�)��	P�]Ey���ы���t��"���N�v��V՟��F�<\T�GH7�/��O�2EH��ty��oM��xF�An��ns�G-k����&,��B%�ua_Y� ���$�;�_�ꁐ�y��#��Tr$��ŧڀx�b�R��;�'pFR�zS�Q)�)T��Ā^;$AA@C�(�eq>�/�𺙣�AAxyt�`��5��]ڑ�E����sz8<a6��}j4V�;��O��ZM+=�Q�/T���*z>��Ȼߟ�6gwX�a�������g x?~8�����Z��6���4�-�4%E��#F3�V��ߠ�"�= ��*Y����h���O�*�L���D�at�������DA�-JW�ݻdv �$A����m:���X9o��a�|s2�C"��_v�cm"v���)�*7��v\��?)�j�H`6O[&���c�3����� ��b�@0* oc@0�8����NЮQ�j�y�&�}r@�l%,�ԃ�1A�z���f�vN,��Q��0K$�u���� �yM�*E�n�O���^���{��	�b1c�z��V��:��:�G˰�B׋^�{��l���WDg6�"�Zv�k�����ŦXa*���� ��9L� K��y�Hs��nT����=�ٌ��ɉ�a`+�{����lc}�X�)Ҏh�&�=��	���<C�'�	Q��VH����pS2q��؋��/ɴ-�=L�����QP�o�7�KZ�W�$��� �S��Zc�H�� u�0���p�V��ڰ(�˱>�_)}�Ԟ��Q�������df�M��@�]�?#_C�(	���=@x@ͱ� k�M]�f���ס�1�_ՠ�q�xm3E�`%�@}1G=ԳN�묦�߾�}�q\2X��;}�����N����rЎjZs�"�:��T�~>S~z~��������m�G� �����m�I'�@#��ћ�m���^�k#�����e��2s�")�V~k9��?��F��=��f����1�����
���W� @ӀL��bD��� ���d��<�kO�#v�O�@���.���tą'����j��[�& y0��\�	:��r�|�"�t
h��D͑����L��:	PR������# pރ�ǂ�:�
nN��V��#G��Q� ��Z#�yM!0zS]�GZ�b�&*Ɇ���(��3�k�Q�a|��'�5�C"�n��<r�jHm�O%3Mճ�96'��`�z�̸�0W.�)N�Z/e�0��p���!��3)�C�bb{
�� dOU��+}O2Y+Y�J����H�]�>���6}c9蓯����5��UW���YmH;��|2j�a�C�X�u42��*��wG�0��c���^���j LmLBZ�0NP��[7Rs�=��K��+�3��F�S�S��&R�P�A���� 'I^�� f�~�W~�<�r�X�[����Ofzw�0�p��u�bW�ՙ�Q~{ܙ��<CɅ��]���j�_{B��D�Kg���v5���D;Y/�o�Bjvtg1��Ҕ���T&a���	��)	�M�`3��3�0�a�69�	�����ں�	��עqӰ��0�g��EC뉨��Qq��D�[�׌]��#���?8-?�0| �ACs�xS��<���o�p*k,��	\�78 �@sRQ���}�}����R%��몢��a'�·t�{�E�,l�eD�E����c����t�r_�G����=s}�53�?�Yl����6�;,���w��O�]yn��f�	e��7o[�m�.�y�]�;b�,[�7�iN���7D?��<�j%c~�G4��5R���`ܕn-���s�%N��)���s)�%��^�"�O!@�p�N�n�&M&�Ff���d��aG*q�y(��EB�GS����ea�u!�FQ��H̵�{Can�������Wٗʛ8y�	.;�&��1�dU�q��^�Ч�zsO���6��7"��4IG�@�wҘG�A��*6VΨ�Q<;�+��9���L�p��Y��|r�/�͜}��h:'�:'�K�!i�|!��Ǌ��J�r�U��5�T/���g|�����$��~��kW�x\b��7&�p~t�'6
�{����z�nsYУ�bRQ:Z������ێ�� ��]0��8ιF�mº�Y_]���$��hԴ�s���8	F(�ݥL|���:�f]�����ޔť��4o|�F�n�IK����c��9���>���g�t�є���x��s{��M҂�lE�;4dz��{��*kO���̂>����>��r2���o�\
z�������kVT�T������ҤZ�-��N$8���-�;at��}���hu{�՝E�}�oaNQLG��-.����XC�rpC���$f�#��n�.Z� @~.�,���~��~C؜!�r��-�I�P�U���Ix9P�ʋ�����g����$WE�M��9*y�X$�V3ǘ��"����I�4��|%��!(t�mb�P�z��!l#Q0�<��[��A��b��~o{)Ҝr�S`��vP��Yp�	F���}U�vP!i̓'Z����b4`��nYi#��>�L���o>�e�
F�H�	��P9�i%�(�=K�@�f4Vw{̲~�3�O&�8��@�?�9.�*J�K���l���L'�;�u��%�G`�|o|�=_���As4�E¸�AH{���jz#���X�>�����4,�J&�7��\��b���ORp��Z٠̔��>�a/�![*�d͎���04�O/�%���|��z�[1]�N���C��j��B��?�I�yA��kොer�C;�F�~��h��c�j1y�xi������C�����z��y�Δ�hK9�}�_�G1G/b|����<�����dҡs���)����*�\S:����'v�4�|���酶p���#�����o}$��装_
 ��ٚy���%��%_6�P�jK]��������7��PK   c�X<��)�  �  /   images/b5e46968-c26e-44e5-9cb6-c624e6f7a7cb.png�Yy<�߿��B*!-b�AeK�l)�ޢi���#k� I�H�D�%$��%e�Bb�Kd��<�N��u��w��w��=���9�|������|�?�+���B�\\\B&G�9#���]�˙}��s�$KS[C��HB������YYw��ES�FG#���;p�Сr��R��N�<��\}  �����_P�������c!�z
ߚ�p/����Uj���.?�s}�""#�^���de?y�\[���|ya���SAEMmݛ��O�/�^V~n�RC�M��q����{�?���ϗ�+=c�*���#���T�@�V�����*A޾\?�� _<�,�,�Lt��ѕ�����z���9�3Ø���=���mB�m	!g	Z.r؃���9
��d�l�����v���/�ڜ�O6ZN��|VWN�熬����>ɏ(����L�`0�Z*�WMg�%��QSE���U�)��j���V�'��#Ǳ���mm`��5�JWΝL��F�U�UH~nhU---4F����A(����A�>��5�	~�d����5ޙ@֕������>����Ax_��
��B������e܅�&z��>dV��םD&������?�g�㉙ٿ����ڟlx��������D�5џ�G ��)�S�W[ߏ�'��lI$�ߩ��퓬����������翈8��'oj�ue5u[ս��4��4�0���ߠf$�����WU[�wPNٸ�����B�v%�y�9!{x�݈h_79�?��O�"�q���K������?�C ���q8*.��������w�>e������A��_�م���[ހD�����.�Oy?���{��z~޹_��x�s��WE���5���U�x���֕#�ʒ��_l���&�N�����̟�J����8Q�

�q�����1H�?���,N3��݇8�?����i_~�>�z_���%�mb�g��#S�p�T2Z��.�(_{��I�|��vs�J@�;.T�]�����zB4��`�S���]E%�cɗD�NE�� ��Α�0 Y)�,�ʞ���1S5�YE�W�L�\��:�[1���f��J&��-�[�=�p����Q����%?�S�l&,�G>,��/�X?�%#&�:+u����%J!�L5��/�S`��}8�L9a���V��u�����A��N����Ð֙ ߝt=B:5�<ɸ����c�'e��|�_~��G��=��Bݓo�ڙ��ߝ�1n� �fN��:8~��)�X�B��(�q@z\���}�;�"�CR��RŖ�M�y�Yka�[�ج���'�[�J��U0ؙ;����{Σ��{��?JL�>��r����rՀ/o#���*U�X϶��Bp򷍇2��m鋛�>���v���j����$P�N����d=��IרB<9j��vQ�a��j<j~�SsM�Dnq?Y�#/ �x�f�VI�#Di�{56����UO:��FC)m�z�;�9�:ή�y� 4%4�f�_�z�Z�[����=��*%�4��'���QCg�'̲fI�ȥQ�)���D"n����|��� �
L(��.Ї6BB"���-���@�-&�o��}6-m,���l�,�N/�I�i-�! zsE3�Fď�P²���:�>�:t��C��'Y��ւ��gWD0;�a��#�U�N��7��;��B���Y1�X���ëY��dS�l�y���GMԓ���_/_�g�B?:lQPІذ���%�Mu��v�����O�۬�|X�,�oz�2~�Zv-�[2�H�c��B\���y�3������mk�ۅ�ջe˒q������\��kL�I�Q-�=0���g8ˬ,���Ѩ���ݙ\��z�=0��|�:ֵ]
�1�����������\kc�����؏҉o�	�o$���z��~O��a�|��4�֬4`n������EqYW�0 `���5[���&)u[E9Vp'�%1���a`5�*ӮxhÞVp$(��+��]FM!+p1(Ͷn��
n'+�JB,[n�tÝ���Bb;ֹ��X_�.@�p�$%{�QD��jY2_Dʜ����n�!T��~�Hnx�l�?�(���S�!W\9�v��lL�)�M�|�R�.ggayc��i��1��rt��(���J���oYX��zϷ�e�(��J�	_���v�����d괥q��RnM:�[���-�x��#�A��������H����3�P�Dq�urL;�]_nMXϵ8v�ʗ���D�V0�M�;��,[��� ��$���w��"�����!o���Wa���X���T��[״�<_�/AW7�a���xbvEއ��I,����5��q��F���=ߤ��/�e��j�FЅ9���`f�u���)|����Z)R�7ľ}��z/n�w�����9C���+���
�]q�˹?�[�m9�m3�R�����y$6�L`��Ȍ�9�%�(*��om����ZOu|�|��&G��+�Wۡ�C_���
{$A����E�z�ƭ���ȍ����2n�X*5 D�퐧f|����}�h?ˀ���\� ��[@;������D�sQt��_N�ի�>�jLQ�_E��Ez_Yh4�¼�2�KcPM�/����F��{��Ϝ�=/B��$%���H��a��Ø]�Eܳ�Y���Z�*�q��9��&�a�@I֞:Q�#e��{�z�lDܴ�a�b�8*��;� F��񦨴�\���RXI�v�s�0�Ҍ���8�޴�5g�05�d�Aؤ�i�u�tl+�P���v�M��+XR,��
v6+��5�q���,[�
%�@��H�l�+���d��eSm���s�G�+�e�!0�y��
�����@h�S#���d@�%8���O��.v��+��\�6\��'�"�D�r��_;H��-�DJ��w}�(�>ly_w<�Q�U���"���h��%�Y(��g.���l�v���K���.8?�2ڠ�g�e�>���9����ح����(��f7���tm�E}�����A�"LN��zPE?HV��Ģ9�h5�u.�d�ٻ����2���v&.ʽ$��q}��L�^BQ�������x�n� �Spc�C�2�=�O�A�kqkW����mg��:�:�f,����`�sx�7�� ������q�Q��HΞu{�6����;��]�Q~
/F}�^M�� ��M|	¸s�j�Eq�RDN�
�-�3
�.��`U�������Hsc��n/�Aj�_	�7eze[F�*��;C�]����<�(���7~� 5ߏ8rl�Z�[�[i�y%�@���y˹M2�кz����4��<���~IJ�s�s􊭥��?��΢�[�8{u��)�μ��6R��"#d7!�_��}��.����β'�㧡�=�r >@�T^��`���D"H#��;2������XW=�O�ମ�A�(K|
T����Yr-P�(�c���*e@����Y�йj��+y������㥯���4l�L�*�ۇ��J�VCQ��5*ԙ��� �߉ꆿEH k���R��q�cs+E�<�j����Uкx�E�i=�"��e[f.�h�))�*���lm�z���ۇ�D�-b0�& ��pf��"_�֓�&1��bX2��U>�����qcc}+4wZ�/+�é�M��-�A��T$t����H�;��%b�s�Эw�G��+b��;�QVS�:W��G��VL���)k��=���F�N��q-���v@^���N	�q���,)@�E�-�w�lA~�%�XϞ��,a
�ڜ��MZ�H��ݫ����k�kdލ64�����O��WN��YfژJ?�z� %&�f���k�8(�F)-C��Be�ҷ�szf)'���qI�Ќ�:0{��r��� C��u���k�L:p�	s-���R�
e�:���P�W�q��F	����۽���ƱFz�pB�ъSH�y1*��Y{ �Dϭ� M��{d6m�����cT�����鱣�wo
uY�Cu9ws�`馠(i�n���Lov��d�~��
�J(�V^R��`#�/&H�5E?t�o�Wf�4EB^��S}��C7�{��d-���!�0�٩���ҠR���>��@�3��'�j��i��é��Kց��(����ӆR'W��{��Y�[�x;��rV�\S?L���q����k&Np�ܒ?�]��y�d��π �?�]���\'	ܐ��I����^�������Il}'S������i��9�8��)��ɬ���SĞ�\+i|��ڳ>L7�	��"	�<�v�q�a&�q�_6of�ѽ�=�B�-*# �K��)[�(��c'�.b�X: ���?:0�~�{Wc�j����ՍQ��5��^��)\f�l��k��}�#�3����Q	[T�:�EH+G
�a­�2���n�<�tIz_ʚ�r���h��pۍ�q^���hE�	����nc��<`�� 3�c������+�/��N�'C�t=���z쁞&
l���9(��ʹ}�8��F�RZ!��ć�'�g�����D�G�e(�pkA�j��a�c��a�%�{,h�rLK�-�������H�v���g�=O���;���{�=oZ<�����}8'gϸSO�?w��l5��S�b�QX�5��M�"\��w�f��ĝ�T��VJ)�	��]�X\\���<U���hrc�5Z��o^��|TL�ͅ!t�@�!�����ђ�W�s"��Z��:,�y��P�c�L?��V�RΎ��˟���J�/�C��[%�;ߡa�����j����N�v��hZH����6�NuTN-v�q�;5z�j��R�V�7S���vx�����k��En؝T��l�&m�_�eT�5���l���x�.�~ki�`PgPO��3�Rc��:u�7���]�r�e�Օ�9��sSt+27�J)[��)��jqܞ����Ѯ����>.X�>-����=V\�"�dʳpB��r�h%w1��Р��E.w\�2��ɰ�+��KTO��#����U�L$���X��T@Ģ�\�'I�7����QOs,�YUS��� =27Y��"L�cM�
`���]�!���ݨ�v���ti�ʒ�n�?D�Z��M��2�2wBt���MY�8�w�pZcUg�{�U�r�j�L}�^���V�H�I��+����Nk�X��K��^)�������j2�;�"�VOᾉ���u�hZݜ<%W�4a���~����%�J�ښ�=��g~n:��v��#�z �e��8��¿컼�qx�[ �v�N,<��9����[|��o����������|*�fԗ���C���B\_�;��g�ִsu�&
ם�5H2)��Rki�>U� �ߡ��'OQ�v7nut֡`���	���.ǧe��ח#���~'^S�Tϐ�S���&T�le5#��;���}������.��zk�<���J��?��O���g,)y^FQݴ�5ڥ������~�F�3	�G��<�ym��&5A���q����G�M7Q�9:�7c4�j�Y/G_�7�1�~]�ܙ/�]O��~��d'��j*��G����oǮJJ����ŮA�¦a{�|�<;�x�������}��<�^����5�['JK$g�n� ��z�Pʏd ��=dd�Kz�&іfi��c�,.Q�匊�@��,�Eh��MGg-�S�b ��ORϺ�x�O!�y蘭�%L��>�PK   �d�X��'��Z  jk  /   images/c2c03d23-e153-4716-8f8a-82529ca6767d.png��uX���>� **���(%�H��t�3t�����]**� C7R�ҝ*�CJא�C��A�|������u�>��{�{��^k��������.  p.�T �x  �ع��7~|W���f�*� ����5�'B @��
�ۆ�G��*t��ߡfd���J����������[��^��9}ޅׯ;	����П���y�0�����-��/�a����5�ҰB� _����w�~yG4��ε��rY�LW*��/:6so�Nh17<'����
�#^����-�!-�27�MU/��O�X��N';��i�9��9�h�٣�^K��I�����!I��s��
��ܹ�/?I���Cz����p�xj�&m�+���W9Bpq!8CN����&P�.�"�xP֣�^�E�A��\�~�C3�F}��#���j=e=��Z�k�?\@��ޭ�zqֿ������g����f<���^?��=����_y�߿���5���$����;2�l��ރ��!)b�9~����+~�}_�y���f���!"Pc�4>��,�+��gD�@[G�%80p=��������r�);;U}m��� FM����_[4هHS^�?���lI�� o���`Rޔ|�Q.{�J�{.���ddd����Gw_F�?zy �� �U�0u#@`���
b"��x��ԡ��jg�߶���x'?�O����������%�w����q��Z�/-�k���"O�u�����x������'篕�������H+��1�Ϥ %��������g[���y'Z:[�?��С'��Mt�<~�}���!qbЏ����Fq�%�� lf Ϫ�>Z��Gܼbk��#JG'��t��`1�Dax�L<R����ȥ��4=uMM�f��w�_�����[	^�_^^^�c``X��444DS�ڿV� ����)�uQ�20�9�\�и��+��'�,?����~u_M=*a�ݻ�m�͇�:͉��L�1��|����D��W�'�+^���,�	��"������<x�')%�O�$\O/�?(H����w�����<��� ����wF[r.�r��Tq�p�;tR�9S����y�)sʪ�L]]];��Xn����x���=�uw5�I&F��e4+�#y���_���'����H�ٜn�E�/h��L$2"�=��I:<x|�$5~NNL�U�2��_U���<�NT�*E7�:xW:�Kkj%Υ�!;IgW=��M$urS�"��=�s	�1�|��`��"K�dI��d$g
����d�G3����>����2-=�TS�))霢>lT-�v�0´���zn��l�����s�D�1je��퓗���rWb(~�|g&Qr���7zm�i���&�~&�qLb(s���Rr��{cu����|Jvs�N�,��ʹ�A�>�u���9+�$�e�#(晊��3�u�u:�v(__��&��S�h �d$R����7&��[��6�"G�{�I(82[f��_ݜu循��7@'Gd���b�
��9��X�b�8&��{��ч|�^M�gӄ��3,/%<���(����ɑY��rE#��)B�3��i!�]�]j<�����0��SDB�1ޓ��q�nO�H�7�:���w�2r@�
�DM%x�Mĉ�ʘ�,LL�7��P)�q/��}Wa���-�5o��X��zv�x0�ke"�z�̝��7Q���TN�����fWα�o%�r�j���]�^=�2Ky0J��g;����%��+u��i�qss�xgl�4@��E=\�%$T��@��q��U*���V����i�k�Q���Q�(���K��~*��8�􃝍��1jA�;'q��0��1�pqjY��x�Ou�D"�YRA!���,6��d#��{���>=<��?�O��[\VJ�rtXb�����!I����r�V���[k��{>�p�ϸoPo	����:P@��]SR�[�}i��-�ߛ�w�����i�$�-��xb|�M�Maa����l�+�$<244y7��g�vՑ=}����u���64��ug�I_֋���\f���}r�v���G,>�?O~v�Y%<"�)���Ć���#� ��4S���rDT����j�����on�7���Al�Ը.���7���c�[\��Fu���Ώ3�J?#yj�%�܆�!r�BO7�U2u���Tχb�^�'�����L��!�tD�фĉ�CT|��n�f �#�������>7ի^c M��Va�7��>���2��y}�E�]�Z��'�u�����S-A9�P�y���]��E޾�7z��;	O�����L=�>"�VuP��sY<�������n͊����x|��a@�
eݰ��!F���'��y,��av�<\�0��犴�t�{|��DC��D��>��p�����G~T7�ό�D��d���6�˲���{����/<���I[��RP��_͢k�_-VV�ś��d9�*�9����T�/��6ۦ��Y^�MB�4魍$��$t�x;��P�{P;�+������L��9�I�Ab�h�o��ձzdܦ)(��©2f�(�����ݾ�P��U��
�;-�9*����J9����aU��¤����a���=�>����X>�e��h%���о�o�|Lu��W�Һ�������i������+�ٰϹ��}��|���ʄ���K�Q#�+����9��0�
��%r��>mZ|��r��|8=j�s�m5e#�BͰ��P����}�����c%�U�?����âb`��ŋQAAT�c�XY�!�t�&.T^�ͯ�
t=ȝ�(�����8e.�l�O�+�<�2�uqݻ���T���rdt�0W�x�@a.DQ�tg8�?l�H����F>��J0B�i�������{	�`�r���|�����]�=������_`o���/;m�e�,��q�ӕoI$-k:�~��A^{�9��P;�}q�IL,m�@��	Gqfĕ�8.!!��f������I#M�PV(n��Ƚ���$K�.��Y[�����R�w�|��sgL���ɒ�̣3�%AQ�F�8�O[FG���(@A4::�l���Û�y��E�G�)ɀ��"_](w�p��Bq�hB��JP���wd����Li�%�`�ɠ�z����*9��������o90ܣ�$�#�C~��?mRHX`�x����E��ϵVbs��O������ɵ7�ఫG�J���5��u_FYy��I�tc�͇���{��~�e�л��:���H���%���5A���L�ҡ���\c�����+�3�����Pmn�b�Q��'h��,�B�,�$�l���sC�!ě�L;5�ы�oB{��&���d�N.**���18x��T�伶�X�8�pX0\(��C��3}vV��݊�6�N^��,�⾠\ܠ?��J��e�l�''��/CY9莝p����) '.3S���27]f��/2vw�G���l�}����=|�nJ�R�z ��a�����d������� ��ۧ�lĎ +;Cs��C ;����� ���u��?Tb<+��8~��|M��'ҧdO��Z��r淭م.�j��ˀ�c��;����I� �O@�^Y]��S$���iz2�emU�o���r[��_�`�X���͟��}���~�ۘu��T^WZ7B߄�1 ���ᛕ��
L���}}k���܁�[��j���.���x�N���m#��� �O��f��\ou����,��Wz%x�	�?���XP��hY�����HNNN��UW�de�N	苾�$H�|�� ��fy,~ޛ'n=E3�\ܹJ<���윶k&I���\_�����c7,���ڤ�����])�Z[�ʗ�I{^�5|�o�Ä��]�a����߿��,��A�U�=��y����w��,�Łÿ����Ԋ< 0�f�[�޾�%�ÿҿr/�@����..�L�J9�����I�Ȥqi{)7�[�����X:~�}���i�k� X®�J�N�_s��/��
��9��Һ��;X��s����9d����zZ�ĝst��g�}�^���yC&�&��WA~��}���K�/^sa�ҩ������
ޡ�i�S�ERj!�#m����SU^�}�L(�2_
̵�f�LN��Ožr{��rڬ	g�j���m)1=��-|��7,l�}�!�k`�d�EZn�v+�-�Nz��&Ӭ'���-=r6m�MzI?޶�3���d5�d�c"P+�6y*�����
��r�Pl�3����V��3�A,�?=���?d� �'^���T2C�� �I�=��JT4�\X�PS��@ox�u����ʠȢD�=>�7���[Z����E���$=}���)�n!�xE�rr`�@j�I���MƠ�W!�%Ko�wf�d���o^�.��6�v��]�M��c���t�.���0�!Kr�7X}G�n���I�$\V%��y7�D4��7:�}�N����8�����B�emթ��~����W6>>�Y�޲#NqZN�n�f�8�UŲ|����� dm**�������'�~7`x/O'��T�ʞ��"��*Yl,�J�y����'W�E�c�G�__�q�vA�J��͸��<�a�0K�'�D9��<����[�A�t�GY_������]������"zgnI��Z��,���'��᠖��}?P�A��]�I5s|X9s^�B���z��$8Ϟ�cuB�G;��ƈ��V��~�N�)�o�HʭStK��_�[Ϸ};���wg��o� w�?8=2�Њ��_�Zg�h�:c���:�ةO��S�ⲏk7���_WW'��$�sxn����ODcm��8�*M�/��i!��C;g�����[=t-��n���;�yi��.0G��tK��J�Jm�S~w��S�����5*��w��{xxȪ��=<T_��	�S��=�tzoGV���%-�P1I;������n�Zq���YX�^�n~@i�ɮ��C�&��k����B��t9��]'���t��ؓG�1�fa����M*�z
x�ν�l���ƭ� \�t�����0�ĳ��1�LN���;����m���S����Щ�|{��gy�ݺu�}�����[6�<=��<&/hAfI�A�������1�[f~��ȥ��'*�ٿ]�>�s�&5.z����[׆>��d�%t�#P���F��g\��������&�L�E!��e�A}�Yh�6�ަK��# �m�b�h��!��L�<5��5�p�n08Y�FFgd|1� ����6t�X�`m�%�z]"��Q�����L�����w@��y�e+M��i����c�m����l���V����'��A�Wh����a-,�Rj.�N�ΐ�m6��5%����v*�Y��i��9MTɫ�Jr�h'uܠ��'���xk4��ߟ�e ��UTT��cp!�m�����л�����λ��|�/�{'��0�]Kw��E��4��xCN 
���$�"J���k�o+�%��344D����z�j#٪��T��F�B�̄�l���ٔ>��|f[���ZE��$�D^g�
C3���g�����������9C�t�����=�u/b&QF�ǌ:�L��s�_)�{�"b�Tp�9qe����^�W�e��Mf�F1'^����w�j�-��F�ڈ�n��CC�%NHś��h����m�Ms���'�A'�|��
�wq� �ρ�ޤ�h���xk5\�+�7(��k>>��29�bډV*�T{�=�t�K�l��G��g����N�ߧ�|Mն6t���xHj �d��}�i}5����-@~{o/=H��e�yD��l��L?T�������'���֩n�bu�Ǭ�E����#p~bx�N���me�"�X�wzq���|VYd��P )�������]"�S��{����r���E�;��0%�����<�a����3<<���q���?��4K���њ��`?���rR����� ���h%�)�sGbr�ǲ��|g ~)���*��zKP�������}����C��ƁBb��	k��$����4O��Y1a���]:T0u��9:����z?��K����2�"�y1����b+�a�,p��(r�u���`�+���%���դ�"]z*}NÁ��a@�����ߏ����a�Mu��r8�f}���4_8��x k��6O,=������g��w��St���+�G�z�|��mU�|��4?�г�; հ�b����/�9�Ai�r�H ��Vx\���x  �SR�

8_���� ��Ϋg����n´%�*R�����>���V�6k��e�h�9*���sY�Ip疂�,	V^b�K�;�냘���:[�'y�ΛB�x1.�7����Pff7�����&?>U# mנ��~I�FU�X��I��Nj���J�}������T��ݽ7 �Wx)D�.Nu������	�)x�q��i�"�5�翠8�&u�O"�QE��N���/��N��\��V���)D$��'Ol�>z�=�{�5�����̧@��r�n4[��es�F��d4���I��vT�>2�F��:��sE#�����2�ѱ1���cȅ����J�)칚[�9vw;�Q����QAII�ˀ�mܙ�5�>�r��R�mR8��i�ĭ�?mͳ0�o}�R��u��A�d��:��oe���(1� "��)&��x���I�z�2�o��^��o8?�� �B�|9��Q�3�&zgk�����I��k����0�ѿ�/��hl�%�a�/�LN�܍��(:n��ԩ8�ii��%Y�>�訣�Ű'l_�?�����;�kv����g�a�v�M�I����[�д��v��N�w�.c�EQ���5���J>�i���d8�� �>*ĨNf�&%�Lʘ�o\Q�Ů=�����sbFY�g�(B�z@���(�Vx{{;o�#�ܑ��Ӗ��v[�WH>�L����t�
�G��βyA8�<n;I��W6��bPs����RFE B{L��Q.{A��&���tU�ȿ�9]ӹ�ײh�!�Kd�B�Z�8�}�:Qԭ��[-\5�HB��L��S^L�jX���Ᵽ��E�c�
>\���I������1ї��]�ɀ�4����é�W�R|����m�7Th�l�C4+��<S�4AC����^,�h{�R����=����^�ׯ��:K��3�	SM
	��Lu���G��wN
�U�M/�u1��f�}?�8��]�_���'�ą+�Z[[������31 
m.˄�!�����Mm
.٬	?0���?Z�".>�v�?&��/aab �F����6��2��{�(��4���L�������i�G�����U��*sN��+��s[{Z�*.>x�ƨ��ʉb$|����'�U���P2~��S!^(��9�r)o�i�y�>ʱ��~}�$G����8F�{t��(�}C�_��j�_�y0Kv��i[��`.��5��h0.iEE��<322��4�̄�4�]%�!�a�=oN�0H�Fd�\�}��J�>z���9� N��f�ɰ~riE��g`8��*`�UK�+�-�Ҧ1jO�Xv������P���Y9�&�Ĩ���+V���~)D���L���� \XV^یk�)��m�����r|~o1��O�3�
|`�u����S<6A���f�Uh/5�o W��wDA���"�l5M�����ƫ��Ƥ�%O�,홹�Y���ܔɆ��Q��nN���0�cڞp�f _`�]R�kC�?E���������N���g��""u��F7��.��n W��_�%ˢ�]UQצc��92�*9��{�OK�`�{P��kA��ۘ&��m��(�5NX`�Z�9��Q�J�u)�J�8?�%����&*V
�)�Y���F� L����"q������J�!Y{K0s�	)���\���]��B emy�{{�Ue0��s���������R 5r�acc@�Ͽʇ�`-���y�Gu��b��l
�M�k5���|��!��cg?��|HA>]<�u����~>doǲ���)+���|�[%Y�_%!i�_����g����z~]]ě�PA9i-A�KAM�
�6q!�?��R���*(t��+)5$�}�'_������o	��k+Y ���5��xw����n����0>g���҉�qM���UM����d.Ȕۿ�Sxd`1��aiD�?��|F�0��Bō��s5�.t_���uO�6���X����y*׵R�3�^�2�v+���	2��#�ΈH<x�`������3�F�T�Y��vM�Kd+z�j���..�}f뱱1(CRa��m�"F����0�v��{r���
��ׯ_���U�<uO�T����!?�9!�J
��������m<8 �H�P5��s�	.�fk(�17����y�B���*/�����/����_R2���b=#�c��Ou�1擳��+:�<K���ռoU�{ J���
렙��؞�Uf�
��db�7��ؽ���7�౶�(�=�y�;cii��6���c���o��M,��Y Y�KxZPJ��;}*�l���	\Ԏ�EF�I�n�2�%5�.��42-Sa4h	lA�_&r*Bc����ٶ]d%�5��ޢ�� �u����v@D����^l�k�	��S��Ol������p�D:B�]����t9�|
����D��Q���|�Ƥ8����q�˼�l͏��*���D)oPu�7��� ��?�J�OL;�χ�}��}���$�YB���rP�1�|����N�z����{^�֝�y��ԥ�ex��D�e�~�q�)H�W� �b�'wnX�8���%r!��q��b�Oj|5�&=�מ4I
iI�`�l��G�v����Y�f� hX�ZW���h���a�$sl���-�x� {�IJ��>6��1�6�=��������,�l�l��~���Ԟ���-U֖Ž�Z����S:�Ż  ��5@�I��Ơ���M���{˗�>u>'≇H��f��ZXX��i**�/���f@YC�ڢC*d�LOo��}D�ف�~�|# ����j�D�D��
㬹�/S��K)K�E�;Pcu�^�m��2�qpuA�_����}����7H���,-cޟ���^��G�I�<�reP�{:Iss��� Լ!ۍ���7x@�:��?�u���!�Λ�U�Nq�W�(,w�K��\�A���P`P˴�u�PK-֑�T����N�f������L����Uۼ�>9�����ZZ8� ��Er$)0�.���lL����QN�� 0 ��W��H���I�y�����'aG����,
��n"
��f6L����'W�444L�JFA�Ez:r~���dv��R4�"Gr{����l�G*=�E�� �a 3��2���ѢA�2�c���;{;r����܅�����r�\���j��g���k�xpB�B��$P�K6�RV�t}��Gp9�p�@���\�7�1�BZ��o��DQ	�����R���w�ܫ����,��IE�V���2ƞ<`�L��vf>����НGVVv4����}"{̪���Fޥ����+�V�ؘ�8Q��m]��/�uف��U�J^�<����q�Т��ձ�@�;:��N�@hx�л+����չ�Z�E���#e�a���YYl�.kU��b�j}i�.0Y�#d��5�׬_I �2a��8��#f�-��/�JDC{���^��ڷ�ڬ*v�:X}���^J%k!{CO��nf�w��Ph� ���Wt�9 XJK+�Xh��)7=��hay�t����HsU99�;m9^r��h!5�W�ٳ^
����yh�^����P+Ԓ ݴ�58�&����N�qB�A:��@�8�hm
U03}N��!��G��a��
I�9XE;�?�m�lJ�%���C�2�u��H�1�Ѡ����U���ig��1�E��ۗҩ��À�Fw7a��)�O;�tnt�]0���h�-%-��0����DM���;^�?n�z�'��˕���.�8����F�I��%�b�����`ּB["-Y�Q��k�l��oj���"q�tAg�K������������e�@���)xĕ4�kJ�Ri� fAA�#�!����x;j���|2sqk�F.��,�"@��V����gl%�!�)+J���)���YQ�Q~~P~�H���E��Ku't	:������1�~��`���zM�Δ�ez�)��dJ��1��}�e�&��F�J�\y]zc8�>�.���U�T�QF�L1�f��Ν��zE�r;kK�A�w"�IQ��N�]�(e��B��Dv�쉃���
?SBR`Ȯ������O���%rῘX�Ϛ@���# ��P?H�(j2'������w2w�*St�HKS����7������40����uvv,K���:�>����؀%�㛮��k?����������W����� i�L��������S��B�o¼ݥ{��ޔ�(=J�w,N1"(.�i�<	�(��u�)E�ߏ�S�90arze�ΚtGӍ�<;u��Qc[2����wv/Z�gff��5mn��棕����\m�Z;�Ԣ�k��;Q�8��_f����m��$HԖ�2��gA��m�QUU"K����#E�ӱxJ!��Q߸r4	|CCâ}�������9IP@�ָ�\��>�����[�yyFq�x{�7N�$��~1 PH����Beܓ;|>I�Fb/w��5���VG�W��
�N��"1�7�r��5�����A������A켷��&,Z[}'���z�C�~�u�r|rrr�KyQw[��2�Jq�|
[q)N�﶐��&�p�t?���EX���������F"������������ %�L^|D��2U[�X�W�dߗ��!2|�V�dE� �.)�]"-�s6�N��������:�˖�J�E|iqOD���u����UҵH���#��O��<���T1�w==�j�JF�3K�<a���]
Jub�R��ޢBq��������PA�TÌ�����W�d�bi�&{D��71��i;l�1	YtZtX�3��6\_k���@ǧ^0��u�x�g@�w�+���l�,��uH��\��ʢ~� �g����Z*h�L��ף�RZ���@BA����_ɻ���w/�dHh����qwY*z��>��-��5�� ��7�S��cbhڑc��ߙ����i�ux���ow4C"�,�}@��l��q#�*�C��7JjGڱT�}����y�sG\/��gYn��?�Q�<<�,V��$����Yf�����H,��\e=�nM#3��JE����A�ޠ)/��a<�y{����H�>���9,����<k��j5�wZ�����0�E�z2 x�.kD�@��bJ!�|SQ.e��Ml�O���� ��oA�:�3l��-�m2����X���TNd0g�Ug:����Z�/_��ܴ�ui:��ى��U�����A G>c׭�*	�ɿ�9a�`�x�>���`��oB���#44(k$n.5�A�x�m���>���%y�S�dgJ�Gcg�<�X�<���'�vM�t��i��6�c%!�ʕ���<9��0���6�����a��"��_9�e�
��]��z��-��������*���
mi�P}�T$ӯ��4wg�V@�/�1�q�N�x0��R����T[�sat���"�uk�~!������y����.S������@P����ҭ p!+��Cm�D�wΕD�n.oR8q��O���D�f`�XP=h{�gcd9-��BCoR���'jj�y(e(N��ǻ���T��V��7��܅�{h�N���{���o�I=����3ח��j���Hz�0T`�ݎ	�������:O�>];��-�2r�|�y�F`�N�AK`?V��_���b{�F�D�/P��zLp@�� ��k=�]̪3OZ:â�$X�D��i�J�Z��'�k�����JU�هn-��0*��ŝ	"���ݛJ$���u�t�qt3˺��@��@�S��/
B�ޙ�lz��$|
h�gό\"��t�?J�ɦ�p��<��>�x����R�o��1h���"�Y�����ȗ;O淆�6W�	��5�g�!<6�S��"~���#`zd�04�\�<���Ƴn�ђ��F�b4���'$Tu�pM�[�&�{�9��h�j&�LEؠh�'`.�.{�Q+�<`��נ۟�d�&vH˗���_�	�A>Z��={O+6(�����B�K�����e��&��w������*��z��Υ���g!1���M�֧H��{"������$q=+� @4b�桚-��]��G`��4V�������f�~���ۦ9�z֊+Q�;!�vY��\�0�4���5�Kj��wq6�ą��c��»���x�_Q�e ���۫����]�9h3@@i+X���.�޶5w�ۚj�)߳��Q5-Up^�Ҭ��ԙHw�M���\A���3�d=�NU�-FbP�����v	U�u^1br�'��`j)��5�;`F/P��F�9������Eb��D����x�u����/Q;�t��б��~t���5l���{����9.� X����-���@ Oihi��σ�_�"���_�#�mi�� 24a}}�N2�dDأ�X9s�Ϩt�	&tb��,F�R8NR8��4�=�t��Y��*�ƀ΢.��s�x�}�H�u��� ]p�l��XfH;3�'���v�Q{��VW̶���u���>�p}�������d�^n��FJ�sXm���1�-6}	��pi��,wfӪ ��� ������L�X�p���ݍ�3t|��Z�vsvOU�A���mv`�ʋ�_/��\�ؗ��A�׊x;��W|�+�5�
Y�6���w{tR�c��F�C�Cϳ�ԗ�AR��B�5+��թ����PsU//��aͽ��6e�3����|��Kq�����+�*�Y`r{�P�♄d�k�ʠ?n����(�7_W�xr�>��woug��?�O/h#|}dP��e!2Aoy��Uo���-�8�gm2���v��]�[fO�F�]�{�H��p�����?��?\'h4�ϧ�&ԕz�]�<��@�x5X�Œ��zjMs���kA|�%�S�N�È|`������y�W�#�A�2L�!�!�����U�~�&�w�:�v(F�n7F�V�4��X��1$�,��T;��(|:���AP`~܍�h��� �����1��0�'�tl�ಚ�.�jS_9���s��f=�Z��M)�I=�et�+O���A	��q	��BB�D��Ĩ��/B�����RV`K�F^<��͙!�ћ+�M����8��7�a�^�-�M�@�vW�V>Պ���?�� �Ե�|��k�ihh�EZ"ﹹ���|����@���r�MWstk��ͨ9c.���q������� g���"�����w>4�0�s�C|m�?8�ݭ�Ru� I�l��*H�6A�6��-�s���B�t������9�U��������:��'Y���N�G:�5w��5rҭp�2C����V3O��;3�2�1�<��.�2�>Ql�.(P�8���+*".n��wF��{f5H.�S۸@WQSp��a�J
�b�bc��f�x�N�w.�n.6�tR&R&������~�,n~�'��}�ꫜs�WǁyZP_?a��4`,1����"�����"yO<��'�8����]j;����[.⎫c�9͢���_�[��P��R9JJ�K]���6*4�!{ů��P�HDVy.SQ�S�K�����)��[<k��l�!~��_�����L&�\�/���Y�H^��X��b̪OzٶQ�� ���"�o�B�ۥB�2�_���������d|�" (����k����V���h�.�ф?�t��i������%y/^�H��<GD�*�jH,3���\<���5�ё���2��U���tt1�.����g�X�Fd^IǙ噭���bZO��M����m�X���\_��W�m;�ۛjTkqz�0�aO���i4��O�P2y�����S�>F�}?��@�ި��c-�P�:�烂��d�z=�:�%��wA6�g��	����tw6�����tYi�����a�~�vg�zu��չT2'���4SW�ؽ����A����8Ȓp�.\(�����:;�̈́��93k��M6��v|�
�i����R,^������#��@t��̓��_�:q����S�mLTK,�f�q(�s^�Аa� )�݊�O��TP����D7���I^�Mq�|Ȕ;���?ޜaө&�[�3������=4�����	���^�9~{Y��{ʹg�[蠌lop�yL ��ddd��
�����iTAt�`Yޞ1�=PΔ��T?ChS!^�L��P ������Z�F&�ɋ�Wv�����\���LjT�6����x3��Ԑ�j�	�C�yG?�:�؝�
�,|�Xp]�B������'�8��B�[U~�~P�7�Ύ�Y��Q���fyP�䕬�3�4����s�q���ƔE�����L�-�5�]������B����fx4�/����C��n)�m�c�tYE��O<Z?�DXd��&Tpܘ��/�fQ���.��o�4�W�Zpy��Ʈޟ�����[�Q��>�ۉꜸD3�jwZd]l�l5b�7~L�L���"X��@W�cuv*jXJ#j�!��Ud�:��>��1qܷo��3[�7oNŊ�f���L�����.h��Pw�.L,�
�o,�����u����h�Y%1?ϩe�vƾ�.\]y>MH�����h�rٝ�l����8c1�;i�攏^G�|/�gI�@D���H^.�%�5�J���9�n�c�}�m�H��q哵'�b˙�cv��NN|g� ������ {O6�rHR@�9M���oR1�r8[R �oy�|���o�ST}��M }j�%5,F�9�s.�d��6�m� ��d���$���#�F=�p^�I0�@�Xn�pM��E��.�5Ipv�l@$��BX�S���F���PB����{4,���#�v�*Ah]�@Y9�M*��o ��@q�+jm�ۿ�f��>��ưN��6��R�D�-P2࢓��](k�ޫc �m���&a�������bCt�p��㺂���ܾV,d}er.��aq'����i�����	�e���
^>w4R�<Q���^q��}Sej�AW �J<��@`�l���a:)de��j0G�F�����t��@z�Рj�v�.�hH��������2:3Sftl�#Ӈ�K׳z�ݗ�>�ғ����ح$��3���Z� }Oâh��XR��ĺ���������m�
y�{���
D����K(G�ǤT��"	C� �*mtk�a��_oG�R����[�~�E���{�[��M��o@�M�x��W�OPR������#kOߛ�dt+>5��Ԓ3ly<�\�;m��ŵCq�CUNXp�@L��P�Y�KF�4fn�|#�'\a�ʾ�7�q:�h��;��������Oq�����DQ�
4��<Ҍ/�]�/��Se3��T��'�J���>z>���i��y�˥'��T���3���J�,d6Z�j9�4����,�C���}�^/>軝4��}�Wu����q5��K���P(�Ԏ"�h�8�T�Ϸ�z�2�t>��=r3�R�^ݺ���n�dmz�#�p)SMC\YY)
�FХ/���:T������]Ϫ��dJnPQ��bW����M�]�@w�ؖ���YOدGc��PJi��̇�8p���� �����`�|��آO}���?4����˗�5-^�\Mb<��D$LV^��ذ�]Z�	O/m]�b9W&蜷f�2;��0>=��e�����:�. XE��#|��$�6X)����|x�M�.E�e�J�_�z�&L��u��i��8� 9���=j7����+pLIFջ��*	5�A�C{��5S�����ːB��yOt����\'�O�b<�虂B@M�����o�K&��vSMh/�t�E����*�ݳ�9��4��U M$5?d6n,���C��4A�e��[|����6�q{v��B�g&drH)�{��9ëG��y�s��|��o��W�9�2�e�T��0(W����ň�~�g���:�^}��
zq���$�?M��D@+���\i�>��j���q��9��Gj	�kȳ�dԱy�(���~�|C�Gճ��yT����q���iWO��iu{�$�����T1M:�s�oՊ~�b�|T���PߋљHs2��L�C�Ә����im����@�z/޺}���gl�UP����6����Dg;�;�b����c����#ɣI��֛|R���aWLɤ �h�I|�y�̱nb���'���7�gr�p�r�O=�����;�Ĥ�����?�siMM�������G?��|�iB��j�K��vǹ��lB��ʌ2m2�(��U�L���Ѥ4��"h|r�~WC>��<������Mw]�8���LiQ����AY�$�E��e��>�)����'�k�	���@g�X[�GW5aa�D� �w��%ߏ,0��X>[��`�k;�Uh�����b�GR(��<Zk�����M����k���h���E`d1.!����M�$�G=d�ތ�3�6�0~|6�B�E�~�!���ȫ�����%E:[R����J_߇�o�i�y/b����z��H���ԇiL�#iО�s�����Ƀ�6w9��z{��@R��'\�3�(���MaF����T�[束�L�mP�J�2r��@�۱WF5|�2:�PN�ǧ>�� ��T�����ށ�Q�6��L#����J$=�=�:4�AAr=f7��߆���EqP�� ۀ��1�9�+�B�S[Up�Th��{�A��-�^#�����j:�-�6'8���@�%����4Ks���5�h1�� H��O��b'���S��H�Mw�Z�:Y��?o1VE�$�)Mm����I��	0����zG�	/�264�1<5�χ����ܸw��h��3�AE.�{�fދ�O�����gS������	�>�`j?��:��䂚7���V7Z�[f'&l`�0���_��w_Ǖ&-����=RAJ�hɍ8��~�֫W���@�gT(ʞG�=7�s$,��c���{�{��)6��`Jxk���\�k��?���	#ǅ<4���:1ઊ�����ҭ�n9�X�� ��BM�|\��Y�i�ƻ��.��ŉ%ga����f�"�8Q���GI	�X�B{*�����Հ������[<���a�ߟ��|ס������[8��3g�x(  ?ڻ��4!�:8��E��b��%c/
-v�b�t	��{8��3þ]��.�30c�8���8¯! >d�OV��x3�Hb�i�"��>O��O�k�.�l Q`Τ�uXS:N�ix����,]'�pM�7��/,�2*��8�<�u���K��A��T1�;c۲��5A�S^�A�-z�0?������k����n�?I���$)c)[	)��]��ݶQ�e0�س+݈%�]ٗE�e(�2�B��4���|2��'|��5�r��9��9��$��~�d�%0�����,d�;��Y�C�(�#]�-{{{'u�BŁ7�R~��̥�8OBq��;�)'1s�ʯ"κ���=�Þ�#{�j/����"��� �Ȱ�{e=tA�>�~���OFJ�u�O#��*.�E���چU�4��"XZRD ����*��!,,�Ąn���wF"Q�Z�[��O5��W��y�)���bLmZ�K�}���C]Uӈ�y��*4]�p@�I�����������C��l�
BRB���Q�ۉ�NTu�%���4 �'6�˷,y�W*jxV�1�@^@�ld�?e�I`H <Em��a@�L�������A�������)�R���[�+��K�W�|y ��Un�xP''���Q	��ɏɋ2�l������3Mz���WFvaa�M����g`+��D�f��� ���<S{����L H{�W�̟�lr��J�G�y��(�/Q���ڋ��,�1���{�� g.a6���|�<ĤO�|%R
6ܧ�&0)���Ei��3���f�N����]�-�7�k;'�7���\\3�I�� G�|��\ww�ի�A�!r�����r �A�eLɉyX>x�(~LDP_�z�-r�gyS�����qT�ެy���@�y���1EK�^[�T���b���B��-�����܉	eɖ�AR�Mx/��5��^�Γ��Q�x���E�=Vc��@���_�(���Nc($�Y��$�pm�G�גb%�8�a��A{�ن��Ŀ���ʒ*�^�P#���ڻ�c�
������}C�jW�R+�V<jeՆ�����8�gX�~�T\��Ouw�%-uu�C�t>�=��^WTYH]�z��y�J���,3孂��5+���F��C$1�h�-����˃0|)JĀx�{��HF�C{ H�s�jUǄr_���_��<���|���!$�߶$L�6��LW{���>:����Y��ڇ��]�񂠿�X��7%��O�=\��E0���[�(+�-�Է�������`F��㋕B	�ܗP���V��1FK����(�ӥ)�����s��Z�|�Og��^��-d�Ή���O�~Z �dTd��냁��k�k7��'�Wz�
�߬��>e�g̽_/t�{,`����� _l�
e��1��&#�`(I6�Q\;h����F��
yA˥�%�\�����:��W;�P�̿n�Yz�{-b�^��[��A�������-�'j��� mI�ow~!!����Otu��ŵ�K�32/,�ɹ�M�΍s�� �Y<��3���&vf!:.z&��y�B	\y�|���NdӤ�����糷{ �q{#v鎰�Y�U6MG >���p����&9��Vr�Z��̷%&-4�'-��o�<�R�j��<�L�o%=��~~�������
��X  �~�M��u��=�<0�&�Y ��� �}Z�Jx�o%j�vy��p<��$���H§��O� >xC�e���̊Y���ᢥ�z�c]�uR2kP��F[����f���3I�U�5�����M�kߑ�46�v��W�£ҡC���t����^��Q�Z�������a��!��p/���G������.��$�������6Y����8��<�Wb�z�>(,hW�^�>��D�t�� 7��!F�W-�<u~m)7�RQ)�F)	�g��������ǧ��9%.�y�!H⪕�8 ���]ڣSW�9?��sf�L�V�U݂V߀�����}�GE�}�ą��џSA£0����@�y����P����I��eM�13a1�gX:�W��$�D�a��%(�������Y�� 8���ů�8@�I��y��Id��r���5\ңlV���NUg}�k��_/�O��l#.	�%�r���|�~���4�z������7#�S��=:���8K�Ȱ�>����\q��������X9^��"�a���62㺬���^h���|����j:X�́K�I��\해��+��Wvb6(y�q�f6ǎ�t��M��)��`M���+��Ɇ6n��o�W���߫%��S�Z[gك/a�!z�[E�㼍�ݘ�j6�Pq[T��l�����w����V��fc�ؔ��r�#U)�l�E-�����
zRL���A2K�G�]*�@J��G�0B�~0�\�o�ʯ������,���R��Y�3dG"�&��t0:�ɵkW�Яퟱ\���:�`<#h�w����K���گ�J�?arY
�ޭ��os{�$�XP=�s/{��#���v�R���!�6����o��6�޿�-�1=J��~�׷BM�����d4!�����$��q����;IO��os�2��1L}�.{C����z{�[y��Dw��D&�'	�Iym>D��{�F�{$"�Q_D<����3�ڤ�:+b�s�ښ1ݟ��[aW�)���:��Pǁ�;mw&�ɶ��u�6��������a��Z����Inm�&�58�)K�>�UO�����O���	�l}z���[G��DMu_GI�����H����!���]����=��-����ՐZn�:����
�y��R�n!�xZ���=ض$�Ӊ)�Z��Ť3�D"I�;w�%�@(�ȕ�_�~�C�u�j�$̧��@�.��ZQ��F��7b���Ɖ��c�EE�
�R��c�2����:���;:���*��4Ǉ��/1��B�9Ќ<��^SSrʂN����\��=.'��u�g��q�}Ev�h�Y�[�Hb�?����i�'�1�块g]u�6?�=�r��6s2�]SF/.e��y�3��Q���(b����t](x:@Gݞ7�����>ئ;�(����*�9�j��w!�2���t���v�[��G)91�i�bĭ����C�Y��?f��Ke_Κ�$�� ���ꚝ)W�G9��lEC'�q�cZ�k�%^-����G>M�~A��9��+�ͩ�5:aaa��@����."��P7�팹%���[���[��[�)Yղ_�HƱ2G�lq�ä\7k<`�+�X���e��4��\�ߓİ?��7G���zc�Cpgd��-~Ŏ��k[������t�gʘ�g?��U�GW=ѱ����$BGw`�h����9!e��/<x0CMp��&Yƚ�x��W��u�_t����y7ūOٜ½!m��N�V���᝝����R�}-�mk�_��m��b`��ج<7�f��.�4o5�z��L��z��
�%�O��ۋo�2�R��&1$F�(������ê��z>R������!l�u�BV��h.n�
xi�]���
�ȝ�>Xs��vG%��F������:��g�g�|�^�Z�)�r�os3p��x֡Y�άCsf|}W���o�i@>`}�;�{��V�U|�ϗa7	7F�O6���{^7##��T�]�Y����*��� ���a 1�ˁ	o�C���m�pt�#*KFl;9z���!^H�۸�<m抃�����+iJO%�h�>{vd���<o̒B�C1�'z����:[���(��<.��љ���e���m%@�9_h�	�4|�2�#�[�n�T.P��k1��3������Y;�?hPn6��O?=��*�+���|�5N4������U����G}��w����>����(��t^򻷷)$b}_�����kwwΦ���m�N���� 97�T9w5k&���Mo���f�,���G'nN���#�D$����5�/�>4��qz��)�������1��d
�9�b��p|%���I�w�g��_�S{@���#��<L��L�<RӐI_�������@�y禚�O���������n�YU[_)
���R-�q�+n�U:+��>��K{�"E�W�~|�5����[5�c~}�����Y��v�N����;��e�%���,����!����`�6�IT�92z}"�měk��T
/A�n���%�. �{����>���w�7��%w���IйF�P���a�l���\RUuu�<��P�����B�1�d�m�b4Mz�	=`�w�|����b�wa3e��O�J{�z_uK�v�S^W�(�\��!z:3�Ͱ�퟼谡w.�f��l&�0a��m����گf��S�):(��rͭ�~�s�����0u_=W�O���Q����+dg��u�Z�q�'�w�W�z�F�Ine�KQ_�z�m����S4��0�!rw�ca�Z�<�l�\*�M�Q�g�����zcSS�,�	*px�|g�	�I������o��!�;��ݍ��;J�(�e�"�Uݱ:�m�Y�CQV��e�'�s�leN�Q�燢���Z��
ұRV��n{�^�f�z�Q�)����iBv��&+�+�;#��/�<���I�������a�o\��S]S9�	ǟ}P'������-]��k}��rmޤ��2?!v�❂71}���� �?J�˲gw���Ld[��!�k����"?��7��Ӫ�	�B/�լ��:.�g���D�,\��s4�,��GIJ�ꕗP(4���T*�s����H�K�r{(x��L��ۂ5�痏�.�B�{�T9/�Qg�p� �ʇ�jߒ�L~�"m�|io��-X��E'c���ё���!`���3,h��O�z��x"/��J��,����0S^Dxx3��7S�I��Ȇ�I�u+l���P���5�7��䷿�Ar�	k�W�9�w?����Iqt�?E�p.�k�q?w"m?T0�_�|�����F�0<����´6�޸��8�5{�)"[yo�?�G;�zx�!���pn�5�ȝ�N�����~���/����"R�O�\� \tϳ�D��EDC�<��X�ݍ��T�y"���ħ׳W��������
���1��Ė���QW)��N���2+�N�*����6N|P(Ă�ډN�u'i1N��[�"d!O3�=_����������*���"��}��1U�cG�f;}]�͸���F��(î�?=�������>�wV�G��ў=�L9v�r[ǁ`�2x»3�j'o��������4����Ki6��ߦ�g߃@d�`D"�f�B�͗�F��l&�+��.׉�����qR��V��f��U���toA{Kgࠀ�ֈ��E��:��{t��y��h=�4�"����I�:�sf�0��)8\��hS���.� ����=�Q�?ͿL����e��%���fJ�h�BɲꚤK�����[� �+�
�n��PK   6d�X�Rr5�  5 /   images/d706f58f-9a00-4cd4-bd85-1d2b1267c556.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   8f�Xjڎ�]#  X#  /   images/f05b9ad5-5094-4ce0-9263-d8ec2a6ced75.pngX#�܉PNG

   IHDR   d   K   �"�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  "�IDATx��}	�UՕ��[uk�F�Yf�5Q#�!1�D�3��L'��tZ��/m��b���D�h̋C��#��"  �XPL5�s�y~���ܪso�*��x�m6�����Ϛ���9X��(�����+Ώ���!Q�2C2�d��/9��&�9^�/��9zd��"s��2�8C������2#�"�����ɣ��PH�1Y���	�3e	�s���9��-t����	3��s�u��Jd~K�?ȴN�BX�=2���95�i����̥g�M!L\��u%�V�v��1�(�(
n�μbD�)_Sb1�rD�o���j���˷$#�0�(��;0��"��'s���2��sj�C2�|Q�9�E*CxP3x�K��@�6�+e�Y��˨(R,>���#�R�P��{�c>��l:C��s�Tb��-C�=B��HL�0Ĝ���{���ʏ��F=�V[��r�+W,Gt�.t�{F�!/�����-}_�����2�&�z��-�׆E�z���`�r�t��_s�f4#�D\��\� Vy8IM�����x,�� �ǰ�,0E"8�a�͘BA�e�
L,�d�e�\�;�E��iO��#-����̯���#C��ts����ΐ��:�����{a]�ͫ�^$=�/�r�����_z�U��-J�@9�$s�uיi�؄p8���1��0S��)���ˬP�L�W5г
����7F�4i7�EڡE_��w�/�L�MRXlQ
+��@�&�U1D=;r��2s�72~�}��h�iE͓xcd#)Q��7n�����oD��D[�`	����G�{��4���}i$3zq� +��IlEZ�Fm�Y���0��	-�R��FN��9L���I>�*����ӏ+'] �:�to�Ob��kO�Τ9�� #.Z�9��ð<G�S��cbry�Q�W�\�7ۅ���}j)b��Y$sj��*�CyW�X#S��ȇ�C��j�u;���IB�q�	CS�'!��Nי���gvdH (����Фl]���lv���G�kd�i����X�d���M��=*�lr0���3HOg��0�P�5�C����iBF6oDЙ#5:2��=�����ED%���(˜IQ�n7BﾅX]�,?j��h�9�_��#R�I�3º&�C㐫�Z�?��;�k�N�����_���$l4�ӿQo])��8[+���(	!C�]p?��0��`� ������i�}���M�lh��Qf��,h��{2/N�A�2~D����2�ɜr��K�=���O2�2����2�v8Os9�2���8f�|Jf 
V@l��9ҍ�<e4�3*���g0k$�M0�3��b
����_~8�9��gH<�b㚪�"q����«�Ű�L����%y�9�����$O�	�!&&�x��Y���	�ǯE=¬X8�^*�,��Ca-h�2�1=���h��k���9�Eb��_E�A�Ǎé;�(�:�O���r�QK���VjE8+��-��LK�[�A���9�TZڒ���9�b6�!X_��K��t"���3�(f��A��UC�­�O}�1�hnh�e�n�#�c����L|�E�d6w����wVJ����E�Y�m߷�U��%?m�z�"j�����"�������~�>t�_�1׭@��o".��9}�=[?@�W���'~�HG�DE6x'LA�|"�r*v��8.���F��ʿ��ezlV�yd&-"������a�f8�[G��E1Y�2�:�]��ƭ� ���p��d\0Q��9�5���������;r��� kn>��-P̳CLѨ���q���q�Pq��*�:�O#C7Y����g0�aĄ�� ,�a�;䐨0xi�K�q�_�11�G����X�;�+�x#f<���6��a]�d�FE�x8�p{B������BAdN��������˱�X,� 2���d	d]��랱�[6^�N����'�6���z��,�� ����)����EF�6�"���c��%BA�)4.�hŜ'V�i�D<��w�Z�X�Jbc��������1��?�k��!c��I}�:�����?xP�/��v���8�>N����00��QiMD�X��wN�������k����CY��.װ.���)�y��k$n�7\Q�������jDu�P�T�В�Dc�_<����$�{+A��3y�����}�f���ܼ�)�����>�|ֻ�#��5Q���G�fÝZ>K��^ɦu��]��z�P�d�Bl1Y>ф��>��h��7^���M㒿E��Y�7s6�gFw������:�=P'2��e�
�k��y"�gb�v˝��f�}��H��r�3%�����!��z�̨���aU�k+�yc�Ӥ4����:��}]�%�B�/��zD����F	���T�]H��!�Q�HT�|� ��ZT\��{�b��(�؛�Qa=��2�,��q���j�)N�>$��Z���+�&MDc瞤f����ȹ����T�鋪`eTFB����s����ɪ�x�Fji�h,�D@v4"Q�ȟNva�3�T����f�	G^9yI�����^���M�r��Y�-�7�N�r�v���S�5o2%c��c�~���O0S�s=p�,�kL0��/��Ջ�Es�5g� D+\m�d�<>MK�s���HO7�"!j��:b�g�0gf�.��1��c"b�'�o�M�?M�?�Ӝ��o�)k�9Ջ�����!61�����\�ʨ���6�B�_�a��Ym��m&~�QƦ�)�gb�� ��7��I��]ϫ�G��D?�IKD*�÷r}��%���8b1�1������膳2�t�F�r��Ë�UBa��n]4M������DV�3&�%?ʙ��F	U��^��+nE��	��jA�A�;�ѻs+�/Z{Y9|G��ϡ��'�k:��#,-�iɕشu+�������3*�=o.Ɨ#�a-��@|�
��.E�>���XB��V�H.��%bd�U�#AtJ���g�s�9u�ܳ�0��g�(te_��:D�݋�;�{��_s��'��@���(�����6=�8b�A8q��ۦ���e(�Y!8�aG��)�_���ϯAVC�.oY�S��B�N�JD�����ފ�
��d�"���4�.Y��_�1����A�of���C8��#X/�0TCE���/�`�4�l� aQX����ٟD��}3ڳ���E��j� BA�Z��'��@-��|�C(����5w�j��n��W��@m��i�О�>D��Jp��xOQ�ʈd5�}_�ߪcw߀ٿy���YSV�9pV�h��N~--�@�� ���;Gr��4;3T]������^R�`c���N�?��{�#���j~��u�m�.�4�)��$�m��M��T�{v�R�}�Fd�@^u��mی̚��lQSH�[�c�Dto~�w܍�7�$��pZ��`3�!���/P���Ҝ��3?(��Z�AAt͜t5��Ǘ<�|S'�Œ!�DV���sT�Y��K�&�tnx=[7a�7���{X!wEv�xzѻ�#dמą�,�GX�S��h!.˭bZ��]����O���-�|�Pox��E�{ɥM�DW��n��]��y��D���?����câ	f��]�U]��ɣC��h�I�	*��.���W�BօM
o��1�ʔ5���{u�\����̈����ya��K��G(;3�fJqOO.����C���r���'��ۜy�dd�B�$����z4?����@������<����-���$cC>�>�UcW����0�2:��A���iE�0h���6��X��X�\���������&�lQK����t���^���k�d��	����o_�Ri�\!�S\� �<PX��h��>#]���U���M�%�����*mZ�Ff��W�ey�D'a-Vk����<f{`+��܆Z���σm�~�0�AAP8��AcǢ��=�q�W���uaȫ�U�l$���􈖛�!��Z�֬���+f����(��{x?<�j�Ek�c�4f���)fD�����9EN�f�Ȉ��Sìi�q��CO�5�X���DǎGM]B�IƮ�ƈ�J�hb��1;1� ��ζ��x6GLB� ø"|;
<��ԓMU<�-dK��������R�����p�>8���ΔT|B�j<
pj�k��2���!�Ԓ�h�@%v�_R@?F]�Ս�=Q����I:^ {�Y���Di	�c�UD�D��\0%�>��~��������P(���� &Ξ����S�U`�e�|�̘��C,��#�gC#�z��}۴9�?��c�Z�%��4ά���Y&$7�%+tQY�c�E�KDa��k~�����"�h�4VeE�?2Z:5��L�gb�o����i���]�'O,�uD�Ø0+��+�;rq^��Rt}�^B�����[6�}�-2�LUX�������v�\����f8�����\X̖�Ȋv�[P$��= ��?US}�;��yc�6u���bNK�:W�����R��do9�,U�A��8����5�B����R��&��ϯ�ykQ�u�e�v�,aF�&f1gwΙR0�-Ȫib�kA�%s� �l=p�/mn|��{�O����̯������1�D� tP��*8'M�M�������!k�B4>��}�o0n�P=�����e3����/�E�&F�s5☴SA���@r�]�l_C}��ƠYʫ;�i��R��u�\g:h	q�	���Q�寢�_���/ᜯ|Iǚ�1�[?@���S��
� �����׷=���\6����o	��[5`�v����ӱ`z��b�$>~�;7���,8%V�>�@O�녯�yˮ�{�N��?���_R��L/�!��&R�SN-z�Z������6�9c�%<p��g��:ۃAe�ɔ��*��:��G�Cr$0�g��,=ф�M���T��C⚖�ΦK7��x�>�v�l��J�._����C��[iK�G�2�G���߹9,�mi/<�C^�z���%�>]�ѡ�W������ｇ	0G�G��@]������"P_�������J�S+�:)��V��3�P�NͰ8r��*rhb�=�MZϯ^�*��޲qIb���U�0���O3Y��l�&�mL��r��ϼ@ׂ�$҆����3�@�CX�VN�]<�n�#MI[�h�t�C���t�2ѐO;ۻ�?Q>�d�!��9�K��ye�\w�aS>�)$/��2����]�m�o��vj�P4�#X���FD�!��((D8�Fr�!&�KN�s�	�t�1i�^�
�jFw���t�аiF��=~2�/�V|��H$��j�
T#:6t䈉b���?�>v��;57)� q��&�MKªRh�2���o���7>C"�WP��!U�U>$���~���@Ԧ e��2,#���^�E�V��$�usJ@D��{�{0gd(�fґ,��y�$���hx���:�fC�`,D�巢`����]����Mg��t�"���S��H��(�,j�<��!ʊ��Έ!L���=�7k�wv�(fֲ��*
��2������!eML��,:�E�cZ�����-}'R�h��d,Wi[^�����Vw�[�,���Vb�8������Ӈ|$8d���1�䞴8d0��e�L}�������O��@w@��� 
���
h��3�$}����r��$QI�FUE#�U��%�3�|�����P�9�d�&��v3T��5̡���9&K����)���Q3UK��X��G�*'6��QXC�:�׬�EBZ�8.�X�#��J{��7�ч�,�8��E��]԰A��Hb��8}���'3�k�[{�����u5�0��*�MW<�N�+��~G�f�G�⫒T"i�ΰ@u�r�ɹ�����/P��;��y&D2�s0#;a�6M@Sz�HhbB��ݪXE��ŕ�>��9*��H����m��z|�܌���*�vN�N�Gf1}'�)���s�D�Hk\�+U�iX�KŜ�ߏ���JjliZ����F�yz��E%�H���dU�NߐeX۔~�h��eX��H� �����=Y��H�s����Ѧ���Lx{[��$~�+��p1�{v���;ᯩRB���˪����]B✋/E�oW�v�A�xa���:��{�2Q����J+3��md|���?�Q�����aV:;�ڏHnLeLV݇��n�V�K"�C��0�m�������
�`4g,PQxx��Z*���@�!t��[^�5ֿ͡����@�Y�mzE��{�mF��7�WExX�#3���*#Nq�c��F^��QN]�h�d�y@�x�?���_�)T��1憛���oQ���UZA�e	�_q;ּ�����)�Z��\q����������������jL#�W���IJE�3�� �0�5RjI��{>�9��.��3b���4�Lї2�e�.����W}Ђ���-��N�ͳ�
z�)�8m����T�gϮ��R�D3X9�X󆪱n��HH|���;��%Y%S��{�G{C�[��h-,��]3�NA����$v`q��Z7m���qQ�a��ab�eK49Lؽ��l��=+{.������b*��ZQ�y��b�e��uo�t嗑s�����"��U+�w����W�Ǆ<�L1a�����c��0<m�;2}����Ȝ6K8�G-L����shB�MjCt�,e2բ��DX
��:����2��g�#��Jbf�:�Z�Z�*��¶d�D�3ON.�z�\�3h��e[��h���Ihwԣ���.>6O��*�x��҄{tEx���Ȫ&2�9ȃ��!�h�Sm>���_���d�pW��Vf�F6��z�P���LGψ��PY~��c�>�MRDi��ogX�9]e��(=���'a|�+��:��a����a,h�JjR���7M{�YE:t��+���P�� �S��A�z�K�M0X�k�o��i:�9�wuz�@9,��ilSE���2�;JJm<��cdC[n(�(����pcb��}����-�#i4R�3(P9<���]���h�3���(����9�j�c�8�k	52����[A�5�1!�DqI�h�|�I��v�.�Ħ�Ch�[����۱�*>d���q`���������krP[��&��-UKx�L��K��?u�ʆsF� �*�V��n�˽�S�����4[}���=r�wߧ
����a��~Au/�Eڻ����
�\q�+w �Z�T�$Ӳ�]�ܙ����_"�۫��2�@U]S]�i�5Fk��DA\+9�hC��=9%����i�kb#��Ť��j**���ke�Y�h]�"&|�G�~�A8Ǝ�M�3�
���������g�(�Uۤ���dL��ޝ��(+WH���k�|�x����E\�8���ŔBA���:�k����*f�Ij8����#{�5��J�DJlA�	�kRT�%����G{C�.�!95����4��툫{,�5���XQx��r�}8D<憛ѽu��s,{��ZϚݎ���V�O�	Ԛ�'�S��Tz�J�v7�e���1tnX�
RL/���|X��VV`̧W�k���Z�P�>�k��[I6t`+�Y��'���uUI��*�\msႬ<X�gDlNS2��8"�����Ml��ǦV�����E׬Q(�˳wܻ�#"��[�<�wkf�P��i0R�{�θQN嗠��j5[*�e�M9l�˜5WB�GJ����|�P��>�l���(\���G[P��۶���W�>�]j����|�-�>YgH��c�&L�3U���-���@()�J�K|V"����w�?�4(Z������L�nД��Ϙ6n�Mmg�(gI��-�C�T���Au0��C'���g!*a1���f��tp�������,�3l���<����Zz�4Ţ�F	����כ�������$�T���*a�1m&:�yK�C�_@	>��?T���e�-�����.�r֍r���3��liR�Gs������l�7��zԥbp�dJ�@��ޡ��R��L��P����Fk�x����x�%;��I��cX�ṛd���Or�#S_w�}vc��������,f��ܜ�xK#"�Q���n�/ �)>�Oσ��
}��G�D�@Z����L��Fs0��N���^x�9�:uJ�V?��o���W�©S�{�gp���c�h��������tb�'23���HnK�$�.��Z�w���S�pX�� U7"@��K.G��I�&������qVOzC����� �T��2��l�a�V�����`Lb�M�*q��!�잗�]����;�B{��k2�k+LJ�S�x�1̫؍r��P�=�h\k_�O��5�X��Q���D9}��jhQ��b�A*C�f�<K������!s;���=�N�U��R�0�SO�f�S5 X�O��b��nh�J��gG�:|U����&>42�1��6�x�����4<{�����0)������$*f���%�4z��ۦ����%���0d�̎ďRG
S�P��1��Yڔx�`F���MFZ�9�'�?*6���CS�MIO�>?��jZ�N|�ӒZă0D{2�YTW)��~��k߇>�Q��*�|�8����#C��W���h�'[o�Yj�C,���U�r�)��d�0B&�pөOK�12�Bhϙ}9�㓭��30���c�A.�hQ����kR��M�bj�����Qԡ4?L�_B{8��1���̭��O�mB˭��<4��7RBD��̿��)����3�����7������C�TI��tH��#���O�й_�1	ڳ��;�f>��� 0zw��\�ARPC%'���8�������(B�}���DԶL��2    IEND�B`�PK   �d�X-��R  �W  /   images/f94c5a85-a3c7-4a52-8d39-8987b87f6a96.png�{�WT_��%D@JB�F:��C��i�.�:�����ch�;��������s-��a�����g?��sU�ep�ɱ ���}� 0 E�>&�I���GY-' �}��A!��z	 �r�^��&��}�̺x���w��<K�JأZ�(�{�+t�'��_U��G��_��P�tt�ιFY?IN}�'�]�HW��z&G�GΦtjj���^'�"��T��~�qLG�I�O�>�ԇ).<rr�֯���2�E?���.�B�2�F僚P��V	@�3d5�$0�u���f��S�Q��a�����%P�����Kն��(�.Ӄ����xLK���҇�����.����M���Ku.I��.�ax�밍�(�;F9ǚ/ `±E�9n"|����g�I�2�h;'�Z�9�)�!�Ug�]�6;uo���#|�UZw�c��>,�f���4��Z�8�����Ϸ�rt�mt䡉ݷs��ݖ���u&Ml�������/Fzq��[[�d8��NMi%$$p5�3�|�o�#=��x������j�ٰﲤ&'�� �G�����̱SS���[��W|E�����e������.\�§kq�qqIJהyޏ�8��Z��a�A���<��������D�P^^=��1:1�T��c� ���L����l�p���G� ���Sd��$��`3���ZNr����rYo��>;�('��8~�;����uv�~o�]*m�Q��n�Q��S����ǔ�:_��7c�()��E�Dՙ��ĭތ?Ǯ���S�wv��޾״�|%�tX�jTR]��q��o�{A5�	�n���-9�@�\�������`�2�o�����ϛ��(@�4�!�L��n�7�q�Q��}+�P~yݴY��c�Y��Dt�n68n�����s����ܿ,��zyҦ�찷[h��y����d7�R�4���4�+:�\Sd��� 6=�XD�����N^I��]#���#�kS(����Y�s��d�\����+�A|-�[IS�dKM������*nK��iN���������t�}��}��y��������w(M�[�]OUas����O�����3Ni�3��v#^^��m�'�6sk5Yhe�Z�l�X=?�{��.� �X"����ǒ�[[�1jq3,e���[��a�
�@K�S�/+N��g��^�s����A�f�`�8�m����)��#B �J!�h�&\ڄ-ɗ>ZL�3bg\Z>��e��'7�Y�\���|�_~�r ���3J�Yz���ۻ�Z���b��#�1��i���c3����?�qg�EyW��ʊ{5�Y�_z���{-3�RF�jk�ׯ��h�/��k�NO��Rn�+��64��́��?���K���;i�'�Z�LyE_�cZ-r�_�I9�v�G���y��79zx̢Ǔ?����mƺ8�O�� ��$��t��^tjj�j_ٷ�����/�i���+$~i�e->��l��9o�Ύ������wᥘ������e2���Q2��A[�J�m��jnT $�����kb��K>��n���&>~���f���]M�@��1���ǳz%��Ǿ!"h�X�Ǳ�:�#������NtXވ���h���֝].(���7HVEo���H�P�MM;A�؈�G#�&i|5�<K�l�.N�8��tr$��>��MSj���G9���:0嚚E�������?G��_�6m��ŏ�0�����sss��n��i��Ś��X�8Km\��P䀰%H2t��p���m5��UTT$�B ��U �w� �|	!9cn>���|�v�p��f�\�N�W^��g�J�?/�D����󴯞l��=��	����0��8�'�ҷ�u+ZX5�ڥ�VF����mמ��"�����fxd��%O�e��z"����P";;�m:�7B�g<�|\7Õ�M �!�����SN~l�Z���m�r���i�ŌkP-�a��t<Z�|�	V�bn2%�s:�0b	g:�����.*�s����0W���r�g��2�[��3J9j�[�
�dQ�I�9�d�����>K��H�?��������$R��TI�*z��"Ŕ�E#������!�X�1����t��e�絴�L��+Iy��j�ԛ;/�M��\BPݰ���S���E?���@�S��g?4��ȅ��Y���67��)"|��F.,Q�l�!S_cs���,��E);�����%�����М�ɗ���YO���h!v}9�������)"�zx�}���=���k�In!��?晜�~��!�l�U�p�H�Q&�:�#�����z�,� �y�t�P�{C�$��U���Y
�\�qn7;����=M*�>܋�Bioa�X^nKT�hgG���M���5 c����hl�w���=\\\�ָ���p�碢�Ȟ�ϫ�Z����'z��}}I��ՃN�^ݥ���*
���;�V��EʖΌc>��q�h���}�|�Š;��	"�M���-2�����\���[�>=F�f��w���F��W>�˕�,+�QE5�ֶ-
��c#-���՛�y��YY9�f�S�� 4[�a65���Z�%s�����{�9ݻ�����i`���K)5�?��)_�)�e�:�.��8�)Žt#�+ �P�^e&<q�ot=;:(�����=��b�h�W� "���퉢8��L ���q&�#��]����a�g�H���a��	��\���N���q#f�K�����J���*\��v�NJJ�qk���M����u ���b���I���e��g�U�ߦ.��6!F������#3=3�!ἵ�ë�&N��`h^��a�q��B��&L�G_����g"3�~u3HM7�m&�<Ɣ̉��jޅQє���Y?��!��wo�El���2���+y���գ��=+��f�%d�no��'~��:��MM>!!!���~��4Q�[Z�~(j#�$�s^�u_swU�Tֳ�گ��x,lm���Gс��+?���Q�Z�ֈИ��}Yhʐb�ǣc�]��3r	 �UQE�7�כ�`�S���Z�.cEړ9ȩ�����	"�*/��P�.���`)�d>�Y�G݃��e���X�"f�e�&y������V��*��.�pÖ3bٮ J[l`%��a>$M��u��G�FV�oL���ޢK�/e�O@�d�cCH��9*��X�X�oi�)b���_��.�#�J01�X��/Pr���(���"�-���S��&N��[�MV��ߟx��~�4��kr�4�m����"2�q�>��4N�L��=��A����%�4T��-+#p��]������bH:�c�slߩn��x�۔�e����v�m����'�֤�����tlFx :d��ܳYΜHEY��h=5Q�	j�?��{Aq�Fw/�b�n�p��S�*B'V�M�$w��k����QxT� �_1���� �z׎-�����dO��-|/lQm0����>H��Y��u~C�3`B��VQ��|V����:Y��[
���m��g�<8�Y��t����^�8��7Z�b~i�o&ۼ����/�NEx��b�hi7���l�Vzm��K������Ѹ_1%��Y�z@Eb�m���9iiiQ�� &_�������g�������m����L �o%��O'1:��a������fj+FC�E��(F邓#Y��0��So	E����ކy��[��G�1#�X��91DCq��p�'gq����9?!�������r{��C�)L�2z&Ly�0��X�'�yp�7i�"�q~'�G�7X��6[�Ԏ}W�>ϥLfP�93g�����IndV��u�MX������I[[3��T����z^"�|w"�M���Ȝ�L�i-ФL��O�ln�0�ўk���}��t��j������j#�7V_y]W���Pˏ�_n=8�# Ϥv�f��(\>c`+f�eih���f���Ţ��9�� S�+�%o"���"-l�f���~dIG���÷���ul��,�  oڥ�3�����;]��c�h����!�V�����E�sT�O�LުR��1�(A �?
��ȁ����9+ ������;�;�(�F }N��!���N)a�ϴ2?�bXf
��旟o6�|`8���ΊS�������œ�t#;�u����4.@�g�c���6}�b��I9 �֏;���sbg�������^���>+z��KZm�ؐE x��
���t�����=0����u����I�_���D�Q�h�I�)�Y`��
k�W��Jx��;}�\�D~D���]�J�$rX_0������0d�|=�Q��_o��������ֳ��=�3�$�.*T��o彮`�����!�ce�I������GӾhi�b������;V�c��t��$�<��q�	z[���w�����S��m��w�i*@:>B��h��NLJ� v�H$�P�Q����u��P�j�0י���ϱ6�ݻ��44mU������P�u�(�H+���SS̀*99y/�j�s^+ℼ�Z�-��'��"!��B:h�*�¾>��Z6a<e;��`z�H-C���fi�(B�σ'CCC��Ɂ{xT�z�u?0:U�o=�J�{{['`G� �P����Y;X���ɪ-`���h �m�& r��'?���-̥h�V�i�ܽ��bv��C��Z_$H����(�:�b�#6FQ�>������X�6�f��=���ݸ��Y�t�С��d֎�U��F,;A�w�	�����Q��O��_q$����0���J�S�5��E�#�Qu�G��m�����`��B�i��Vշ�4�:���xe��>�pK�LWY��?߾-�O�'��_�/�)|%�����y-�f��E�R֦/q't�E�t?��y`�sq�)������~鴴[�nr[in��i�^�f|*�;�h3k!�AO��f��S�_[��CW�D`��scF��K�a.�f9:U�N�cя>v�������G��B��^�)HI���~���%ƨ+-�弢�,^\�#���Q�X0�q�1�g�ĹJ%��!@�aF��L�P/��%�n11�&�ʃ�"���$�x��`������S�"&fWP,�K�4S��7M�߅c ,z`{���,K�~�� �m�|K��e�Я����Fgz��S���3��&jQ`��\��V77�٤�����Xmr���೗��s����97W�\���+��W�SV�݂]w6��Y/���H�*An���AQQ�>KqT����	�?ssZy�Y��L��x�%I�.��a(@��?�J�X�X'�H�"FLXxEoʱ��!Cծ�ߗf,��h�&��c��H��A@���- ;~��9�ݤ��$T�o��e C �VRFADۇ�:〯��ȃX��0 x������Sy7�kKˈ�C��_��es���r�/--�W9ۼ���V�YxD��'�z���_)�P��'���t�~�>���n����wBHӭ������A��kaY.t�y�dmn��� ��po��x�����~�It@����ݽ��Ç8;]��	\�����a�$k�ʬ���Pؘ*j`I|�C�y��QPq���\X���y����R�Ȩ�Q���L�ɰ��YQ�Ҭ��
ؑ �^l���C��>�"����ao9;���tWj7��3��)�0u��o���X����L3��_4��3|gq���3P\\Y�OFI�Q�M�E?!c��qZ0<G�1|�����(O�0�y���9.;�C&X�-d�x����D����B�n�f�,9R
>��"�r��V^�j[���h��lӽS�oo����
�t� ������Tb�X,����j<�H+B����
���	]﹯�q]d�i����({���l�RI%�oy�FI�Ɣ�e\wqPI�k�&���( ů���&�����xbؒ*���z�ڒ�A��d.
��v�ʜk�W�Y�s�P	�7�lF-� ��#ɥk����+�g��7��*���
|��P�������׿[JIA�KF>?/<���i��1|_Z��Dwu�5����i���\��Ri��1�#x�[�㺕�D9���{��4���,��w�H������^�#��!^�h�I?� c�0j�tB�G�;PDa"������Ői%]Ƒ���cÖ��ǽS���o6a��@L%��	'4,b&�_;v������aaoO¨b�b8%,,���J)hH�v<�&N'{�fj�VV�gߨ�4ա��UL��3���@�...�}t:�@Y���b�_>�{����4�ڹ�ٴ.z�q�E���G  � 5"]k�<2@�l��0��"#�6��h����T�4�ez�w�9ᄺ���ٝ�ר`]u{n�,��
��l ��~(5E�+?��y�J��M��^���@^�0�)5�9:B��gC�O��I+�8�@��p�mN�娤�:�,�y� s���UaT1��gW}�X`J�UK���B�Xad}��?�x9�e���'2l�T��F�T���Nr�m��~9.{шl�� ��L�rt���h���ٙ ��nռ�L/ٙ���œ(y�����������"C��t:������6���Y��"\���}��J`�������X��0dJ���U��I|��xOlpk9�I��ڭu�F����-UΘ��,��Xܻ:wz�UR#]m^~L�8t�]z�++�dp����	�/��u��}~�V���{m�D�y���([M9,�B�I����8I��=Sʾ��oAxǥC퀂�g �^�ֶq�٨�,/�"ŤH=�:��ᡃ
�]�(,�xk,M	���� c���i�y1�tfQ�A�f6s�%x�~���a�L*Hi�A27�DX��݇+<��.KG%򾻢����ɢ�Yiq��"�WK_�uS��D�
���!Y,De���k�j�/�Y��:����Y㙓Ò���yBA�bw��˷���H?���jNQA���]��δJ[o{�#�&�|$��~�����]��+��¦$�������TS�\q���>�_sH��6I��Q�x�ke�H��L��ʦa�fj!����O�����j-�az�����P�o���!�E��a�����:>Fe_T���+%�X=R�.2
OK�Ӣ���t�V��N㇞��(%ҾK�i��6��l(Mʇ�u��='�+	4zo����M�+�Gq����U��sY�A�DbuK�/d��<_��K�mCJ��Y�95��V�rhh�����(,A�����/�Oр���]rV��B�g5�;L�=e#k��y�_����Ix]D��^>&���c'�?��w�b�*�yH�����[��|��)Of`����V~֣,�f[صxÀu�Xn)V��v(\��Ӻ�(�ס@u"��;7������ˏ�!�@����ؗ��xN^.�M��Ʌe���$T��tD�L`T@���BR��i���x_�/Q�nF��M�
B'�"sO�=>��9��	�`��ki!;����t��|�	��J�FG�� ���VZZZ#��pOET��߂؂�R�Q�ɯvR���&�(�m��6�O�Hf;�X��j�m�u᯳�8��� ��	�8��%�`����PS/���7�{�Kw��Odwh�#��\�����:_[U�������2�I��*�,�%��N�k�Np��Q��K�h8��&D{��l�v�T҈��楰�w'h��*q`�e�4�~Ճ�U��Ͷ�	�E1/�s�/�c
+y���̓b|\�I�n�G���W5]Q��,gC�B���ݗ��9��j�b^�������^�����e��W*U�5$V� �������q(^ໝ���佽�Iq�C������/�#��U�0�9����O����qN��M���R�hb?$ה��Ĭ':��p��c@�>9Y���CgW#g�v���{݅��+����~/Ɵ�L�l��/���ʮ�̢ǋ�x��;�����y��Nya�n%+�0���~�>(�k�����u��cs��hG��� ��߽d]�f���w�MY:;_/Dl�Џ0�._����ksrr���@K�u��#/���l����\P�ǐ��Ayٕo��k���ζ�P�������&v^��RXO|�r��ް�k/R�@� `��W��H�i[:�#CH�X!m���a	�����Y�"���JԿ����( S�������B��ץR��{~�$I�����ё���UX�<	!�ňM��P�<iR��1�7�-�{�w[=xA/ȧ�wÎ���G�m�N���c����]�k11�C
����s��Q���з`<]OD���N�+N)K?l�`�"7}ٰp� �����=�_�p���~�!��!���@�B�Y?/�
\��2�Һ|�F��{��aW���|�4+Z�~��|��FZ������J�5��\H ʁ ܇�V���$+�`}yA5��� ���bDB��%S�zb[��'�����4k=�'ܵz�i��dߙ����������i�e_�D�hM�ב��g�T���ͯ--�b�/�vdD8>�RQ"<j8����by
��~��VŨ�p��:ݚ�~���{VS��q=�J��JDH�$Ы�R�Q��5�g�Oi�s�՝��l��sӃ�]��2o�����
�G�)�,[�[-����ï�2:~�f*�C�����n��B�XG�ʺMB\Z 8[�_!�D�����		��H>io��&"Ǖ��u �D��	
05�]���$9u�8	N_'eK������k��Ǡ
���U��I�0��Ų(-��{��:����|ۗ���@��1\l�@�����:���<:U'�ס��F%�_���� �O�`�Uw��+s\�QR}OrT��'��DE�!0���J�#8�ȹ�4�hТH���EK��k<�z��v�&���߳?m"�]�|S��L���˸�y�� yh����8>L䴓Ri �Ԕ3�s5��ا%��8�l*{��Y�++���Z���y�J�}���(ݘ��\��f�+0I�]O@��ih�?�8{������}���3k参��>�pe}x~��"��#IsR`R�y?�(8��� �?۝���T�I�E���Y̑�v��E�_���	�/N
R���~<p ��#���=��-��Z�	$e�z���T8yXPUK��{�#��a=�)�o}�h\�\�������Ȉ�x�g� O9ٴ�gk�o��Kp��&�z�6&��������R"����y�W�g��)���B��2��r��j��6���yZ=�O���Ql����8!��o�;�ⶡɝ����}������
���X�+����5#�q>9 �P0��ݢ�� 
��x�����բ�ˢ�<�V����cT���'�\{VY:'�p��rg<����pG�6}���%�M*��_E�&����;���&h7z�{,�}��^^Xh�Y��L��`|��6�q!2�)'�08���8%^@��%�[��p!��_׻��y�5�_��N�'''�%�R�h#�I��1;����U������a[���j������J��O��_4��Eu�v@��<ݶ�Ǹ�Ck��U�=�G�b�P���I�\�]��q\�٧v*�`���Cx�QJ���n�`���r�����:������?��������}����;�������&-5!!��c�	����Ư����<�,�vجcp�}�\��b�2�Qd��:���m�:g4±�_?=�5W뒄��]Ԩ_i��o�~����?�'�))��>{/��F;6�(�4��hltT��Z���h�N��E �W���8t�z��j�>
�n�K�D|ۙ*�v��-�ɮ<ob�g� �M~��I�{ @�H��ݶ�/���-����7"�7<�ޟRj܁�g�U�w�DB?��' ����G.�5~&Sq�Q
�l�_gT�L�0&	����z��T�!�Pun�7����Oj����.b|:��J޴���x(~]<�c�2^�Ǫ�������[O�8����&�˄Qp�bt��4b����Yi���LJ
d�XG�� ��'��]���YڭF\����V����k�p���r�ĊLB,g "�e�o�,��4s���N7[�x�����X2�_�"[��5N񤸏&��?��0����|n*q�}w��!y{H}���N9A
�dnn����4q{oO��|���h�m7-��|_� ��(�� �~��-}ʲ��"�w��w�^�ԝ��yր���lD�	�╒ӈ�X�{����R&�`$"@暎(U\b"9
0</>�׿p�c.Κv�k�2e����=*K���=���ԍl��(����8jhL|jvpq�MMLM1#ێ����{�N�t�����1�"d_Q��pU�7\��4���i=p�╠���=�u�;�z��SP������Z[�1��_��B�uQA������o�?p�ZZT/}�_d��OT���Ϭ����Qg�2&
��Jɕ�Ny�Q�^��=�<4�������bi ��߼C�Af9�=Ri��]��z�F.J�@�RF����6ϭQf�`K++��%P:kK�R�vvv'J�sK�[kG�9����5h9��}p�����J������b�ۮ�Ɨ�����|�/�u�#�_��ߎ�o1��^qR�7�3-� '
#M�H!�F_J��㼅�?K|�g@���r�h%��zU�E>�J_CԸ���u׸]YR2�o>���sZ����}Q/ �O'���	��]~5�uRk����(1f���G�o��}r�P*N"*���K750�N:9#̀�*r�B��(��AKZT���,	a�U�8�E����q��/�Y8芠�0�����H���ʳ/]��u�Ԝ�7�7�NJ{V	�_�����$(X�A����X�K��Q�I\�>����4�¼2**��V�S�w��� n�+�D.Rr����ٛ������A�/�)%#�ph����7^Z2j���b��9�X�{����kB�E�?ڔe!S3>9��2,玿�I�'c��Û�����>����������m�������gZ��T��vU}e�G6㇓!tK���1��m�_f�#�ȭd�#���t��u�A^w
�']��۞Y����O[�?+��$��V[�If���y�+���C�^�e���)�J�i��+6rG�o)
��mk/~�i���bh���v!uu�ϙ�{��K�"��y����`a$�π���u�ea�Ze(ɍrdF}&v����C��**�+��\Y�:'�Q��L置v��vC����5m�l��,�j����
F��>�!��U�˼k�pN�Ƅ�诓�X�H���aiC��w����8^�q�jg֢ �*RJ���9+�)"JZ��3�ލ	��<a)�v�Q�,��̽y��!<�������h�qy�q.��Q���瓝2��n_ǩ�y�[�e�}F䤲����)����/��(?9���n7U���cC�����P�eI`޵��!�0�r��:`8V�ר"V��3�-`� )�'�U��]�]Ip�:]݋�ϟ�۪����r���,�(}�X�|��D��J2^�n�4V��$��<�j�����Ґ- Y:0���S!��.3�M�o�d�M�=�Q��E������0�;��n�?��PM�\aF��3H5�hn��k��H���Iv(Mα�u��wv��sxފ�#q���ebt4Z�h ;�Y�Ͽk:Tq����<���F|]Ղ��?����(��lY�6������� .��>ra��Euٮ���[\rrrR���cW�V���'>y\�X>%ϯ��٧�9e;RR�cMh���G&ق�[mmmQ�PGR>�XҨ�ԋ������]��J�q����1w��i��M߆�O��XOϓ�w��&��eʬ1�Kvj�FI���K�eL��OEA���5us[�,Bl�ֽ���,c�j��n�׾��3J.�s�.
e9ZO�N�H���O�P(52�(;@���+:n+�X)*�Ȱ��x��T=?r��r��U OA��d}�`��U�ȝcW��@����œO��WJ��ǻK��󳊊
P<�[=+�T|-#�^~Z;�˄0q�:��7�|X�8��^�dd��s���F�XB�B����������h��1��76yS�i�:�?��\\\$t:Y��P��7�������EA��AHJݚ�|Ʋ8��������0��-�_�����^/�;{)N���1`��؎֨�>�X�ڴ��c05�jnY�Vu�.����b4������&#�O���!�����*���"�(�N�Φn($�|n|!&=�G+���¨��C)4$�se�gu>J��i���H�Zn4�;WI�� G�t�=� h*���"W�(��c-x��_���4��*~�z�b>�P%�����!��X�zrh`=��w��T0f��?1�\K��ޱ�
�O���T�ud��uoB�<��I�>сڏ���
�pO7n
S�F.n7�IN�_�ᬑX��M��dg3�]�!&'�vͿ[+ ���qF��Wg=�� ,}yE��0��mv���QZ�jc�b��!F��ȑM"@������a��9�����4�G��Rf��B�|*=R�\kj���뿚�ff�!]��=�^�nvS��8>[<Oº�ݤ���Ep��-���g���WhF�AqÔ�&%�x۟ϭ��i��s�2��"ʫi]�|Z��	�߾�j��k:��%�����Q�o�L笴�a^�5^�t	W��(���K��v�-���;����׮�^"9%h�/b���O3���"w��m�~��i�wQW��xP�����\R����תҲ�K�x;�9Ϳ���Ҩ*���w������YQ����R�ޥu��.Զ���ohV���yM������piҾ����Pܥ����X,��w�E[oE<��R�=�`yZ�]L�8�[���5�X���7��ט5�R�BZ\E|��o.vV��{	�ڰA�okt|��i�yk�z�7�o�-m]-Oް�Z}4�r=����5X`�Js��?^��_ K��^Cr	�Yh�!��D�����UwTb��;������ٷ�=조΀iq�}�O����uh�}��	�H?��� 7��Juc�-g���[�ߚF	_]������,-���<�T_�O���AH������X��00q�B$���g�{#SNE��u�X{�Q6�a�Q���з}��TO>��+�Ź�v��f( 4EbM����bd�2�@���c��k]'�'�\�=e�߱D%n?o:w�_u�9���\ótb�F����-�a}�x��������S�]і��K9��~��C@�5Z�ޞ
@4�����Ij׌[��=���d�;2�1��aä��B����6N�m�<�s��ؤ\qeۨ��=C�9��B��n~���X?�\�Q��=���Lw�G�G9�Z�?���A�{��<=��K�k�!����Z�Z��wKsz5g��U�s�駫(b�o�|�3��6��r��w��q�}�<S<ʄ�9���7�[�����r��\#�  �̑aJ/�	i[f_Ù�Ah���;g���}m�q�e��{��M.Q5ء<^��ҲÚ��8/�7?�|�+j�A;��x)*�~*l�9��Ox͏6$xͩ-��{M�}S�Df}Ys)>�]
.�[���ЀV �>�>O��v�M{���e:�yyzz��dz���8��cgӻG�}qw���=��)�"$T�o[biSw��z(n׽}Ѝ����t�8�57������|5��m�k*��&��P�E�Bc�1f2�6,^�t��ǶD���[J��	����Y8����J��10�����#E�'���g^�X�3q>��|���տ8���j�A�:k[��7�Hų���'�BJ�����۫��BKE�gN��ׯ_��̔JV&�G�Y%%'��*�0��l�[)����Z�Ȯ=_
����"����'�v�<m�V�;�����' �3�;$�e�,vY��
<""�`���`6;��k!���j���h�$��.k���lU��%�窲�Vz�ж_x�Ϭ|��
B.�B�+�˿�,���K�]��r��?zh�ڞ/����{@y(K/o�0�h�U��/_���rI�3�T�k��0iL���'xrH�p���-$�\� ��"S�����|sC�t`��s>��}P�~S��T�s>�T�Xqg�`� �|f��s�S"�����$R1��È�ƙ�y3@� ,���}IX��%D$FÒ"�أYTth�#���o�T��@����Yff���<�<"Ԛ�*[̫cU�Ib��d�{%-�ܽ	B���E�V&+R)+g��`9�D����wv��B�8��!|<�!��R6���Ī	D��t����;�X��P|�s$����p��>��쁉ʼ�]�2�D�>qU��:!�'N�rp»Tdd���( ��ȷ�����=5���ƹs����Ѿ����%Y`�lN����q�(� &O�Rb�cžU��86 #w�Yʓ����E���?�����PB����n�@�e��7����jII�J��=V/:�U٥o���w��S0��2��� ��|N!��c ���M�߲Yo�x�*�'���µ/���-���*y��^3#ո��R=�h�"���`{fǟQ������JQjӱ��Mrrܗ���t�?u� ��`&\k����9O���F�4ռ�,Wf~���t>�gU4�o>$ &,DX����UR��u*��p�Eu�L?�e�սZ_Q�U�2tTM�����)���jx,+L�鮔��<s�d�7�z�"�$��KR����㿃��Ǌ$�5�c@��Z֧�λ�g�I����zt�WG�^�՘/!��Cu얣K߭�I�}���"�|���O�O��W70��S �S��i�si:��M��H�n�9�=���ǟ��P!�"�.�r��<�eC�@i��%�? sK�ӿ�{T�I#y�����~˴�T��8��k��� S�R�R��@1��j!ٯ��7Rf,m���]�
��:P�d�G�vv~#z���
��~�C]�[?��kNR�1=6��+�X�:�:R_a�d��ݱ�����zw��2w���0������Ⓜ\_��:�ÃG���1�şo�_����W��o��Ec�����s��G�d��0R���.2*��0�}�)��BН�0r���8����r�C��ʋ��{i�u`� �0����e��l��	w|2�Ic�B�ޯ��Z��54M�T���n����>l	/N����C��}����ն�`�q�匕�교�]0cs�r���u)�E�nfV���N�j���< ���> ��r�!�'l�jbJ�԰��O����4
qtͷ8K�}�^���`���pW�� bq�X�ث7z�GSF=^��@|�P5Dp�&��<<y{�"@"����(�E�[{܏�^�z�4b����j�/���,�L,�=�g�P�ɿ�OHnjcZ�����~�r�����1Q|�	���|(r]���3��(��Aر:a�S6d���� !��%硜Ԗ7bb�S�ÿ�O�����DX��. �O:�(�lg*;����5)Sd��ih�Q�U�rs�&�)=���o��T�^<?���AqH���o��?����	��E%U�)�8,@=H-G�q��u��ߙ�|!_�L�թ�2���$�\���>�9�{��F�O<��w�'噈"GrT44� ��$8�P��]bK�dۂؔ
�K�r�����|�ӵH��\�r�S�K�jÌ�w�H3a�9ߗk�hL����@[�^�F!��E�@�V=g�>�^��tj�H�ȗ`����ض�mP`�W�r�8����  �l�|cno�/<P�UPq,�$H�DZ�!�lQd�e�U:`���������ݰ�����Atlq�;{{�S�k�yԉ��Jz>�e_�aCi��X�HW�*��'C�e�Iاu��pZ'���7��r���o*(ʦb��6����������۹�K�C��J^CDR�4��>�A�C�L�!�@5�3��9T�-�v
�7�m�6/8�q7�7�עS�5Nq������r[]��>(�L�Pd��|�E�o���V�@NFQ�:i�~E b���������!�]�e��R�.������0��O�]�pm42@�32Z�� ;�hkk�;,x=�2tQ]�UQ��fi\���V�6p�!��C��\�,�F�糫���c�cC�PJ����(>FHT���Pv���E���� <Jn�q��*�a��d��5>r�1�$tYZG�.�ǈ7b�+�q-<��z�s�����9���z�L�hК�?r�"�<��mJBu*m��A
�P��F��)l�ApS֟��:bw[���'�t�.��IW������ƙR��F�&�J��vE}?$ �)Iƥ0�t`v|�����z�a?��VDt�8�8欔�+�+��(E#�{��A[��E��a��NB�ʛ���w��.I[��	ۻ{Б� ���7���o*m��f�n�QT���,���cl��夭�����k�O��A;��<���V������K���깎�2��9�KI��p����,:�u��U���>E��UD��׶���˾17�ta���a�6�������Kx֏`B��������v�0�ڼ����1�:��s9�x ��h����|�neD�9�w�Q�v)�;ln���p@p���Rq��;E��w�M�W{O�?S��:�{�.���¶	�PrMj�{��h��Y!���I��S����O q�M���8�`�6�|��m�4�#4���*������̿�~�?���>�%I�V$��ɾF��0ƾ�=�,#{��QY'oa"c��I�$C�13��m��c�f|��}����9�u�}�s������)wA�Z�r���s�vBKۻS���W����e��PV�9���%{<s�1�vz_q���6rx�
in�r�L>W$� ������.]7�H�\k[[�\~ș�WL�����T��+y�"C�o�Λ��Z?=�w�NF�ƿ@WDZ�������g�
&���8'����$��Ejҹ���qC�GeFTUUU2����'�H�ʜb�m-y/&�����12����T!n���<b��N���S�i6����Z"�_���m�Jl"Ts
�67��\������b����$��(�};q�AHC���F_��!�!zX���M!����Ȝa!<�e�͔<yf����OTg��v��=sW��me�] m�Ļ�_73�;7|^�	)���J��S�W�]�}:Dt��g���a�3��|1����+V�p�%W�ys�\~
�w!����<��_���7��ϒġ���cnbnR���ӗƲ�/+��C��z�މ��+rE��:�[�����|��)[ۓ����'^�I��~�=d�mU}hW���VP�Bt3��0Mi<�q"Up'�����1t2��c���݃���9_5�7Mjov�z5<�ꆝ=YRX��Ɍ�!�������y��b"][n����1͗��ˎ,hHJ�,��.�y�c��5�&�Dܹ61z�SvȄ���=+|�=J2!I3<��;�0EQ��`�î!u�9nH�Y�`9� �;���ݽ�FF�o6�'i \0P7{&W��j��`Mmb�(�0]>�N��^�D��0����(-��0JQ� ��!���bA[-���r�gʷ���uI��[%�;>>�>uu`�7��T��n��T1�qE1K�B`�訣�O��;���;�w������t7d�ReYQ�i�+�Éx�-CWz�R�D"�._��|�u#�\vi�v=0n��r��q�yUkS+�T�<e���m�jה��N\7�G�Wr�"�+lvwc�z���@hI��2B�f��nvf|'l
��RNovpҫ�9'�1T3���u��Cu�d��x��|�/�����������Ʌ"t��<�Jmni����I��{˳��� �;:z�iiu���0���֬	�[��W"5���:�^�����\��tr��Pj�ֳ��Tһm%j5�
�u��w����Ѭ��QS���_��<��.Q}�X�=�?�����V��[���.pw�d����(��j=�9�~���"ޭTF��)ӯn?n��Yo+�_�fC�_����g�����no���C���Y?��˳��A�*l���6M��8�2�1Ά�b1�#OT��]�x	�uj��'�E*g�(tsx=/�()�$>�g���*���ֶ&��'3߯�^��g/���!�9�q��M�nS��cC�8��n
�&�ѕ��F!w�1w�h�P�?�{���|���h����z��T~�$` �V�Q�1~`��@�Ԓ���d����au��.}�4���_�����P�Ԉ#_�ݸ��N�Ʈx��Q��(�����g��1	���d�s}�i̧3l|ڷgn�S�hV��GN��e��/�ߠV�&d��6��[�4wB��<2Ӽ���'��,�oN�z6�Q���`��us������t猟c�a/T�~Ze�� K�p��uLͥ�[C����������$���ř�>k�e�]��ˮy���}�c��|؂��n��װ�Y6ׇ4�Һ��� WB3�B���A�Ѥ�޵���D.?��|:�� �pq��g|�/�D�1�>�6;O�]��X���=�T0
q,`.������;�C���-Q��Y�i7��������[K�a�����<�f��t�s�Y|@�D2���\��>�u�D`\WG�B ed���l��BD��3�ie*fR¤N��SMKO���^Į9�Ig�y��XlK�ωv���#@乡�;����>\@q��W_����'�ʗ�nG�j����]�<�:�v�k�Lݗ�	p�5hl���̆h2�'Kq�LK��|������&nQ�K )
5hmh�\\\����o�B^d��E��ޟx:0�(m/<�����
)�\if2q�ћd��ٯu0+KۦK�#�ڠ�m®SKaE�Z����\�y&ތ��D\u�ǡ�? �?�Fomb ��6!_�A����o�p꫓�h�����GfJ3�c>���̼Nt-�i'=��l�.U3�݁��P�
}��:���Xi���ߤ����)>iH|��ˠ.�S��e���Yu���&�F�� c����e���N PW
�UPP���϶����Yݟ�wٳNǆ��Z��Ǩm�=����̛A��mfM�q�������kjjzNEFBBX�̜��4������~��v�x���F���>��j�/����N���v0Ƽֶ��9��P�B$E0�7��g�n4��Ţn7G���> '5����]�N�xf�ac{��z4��3�����B"6|�3��$~R���#����km�%�R#�R�| *7ܲ�yƱ����^yy���v;�7`P����x%��.�Y��/⇾0`D�-	@�Y�7��7�/١M��D7���=�N�;%,;�q�wM�8��!;Q�
�oߦ�Yz�!%!*�IGR���\��;}	����*�2����m33�~He�Jc##O��0���
�B��z�r�6��/:]��V�+pB:tH�M�0�ԭ.��j/����!���z��.n�m���P� �����p`���IIK-EOKI'��f	e�y���'̢����>>�n������G�Ɲ{��%���;ϻ��k8�Z_��
2G��ddN �1g�q��.�ASLDXH��`�ڽ�����tw�;����Ը��d�X{������VDaƈ�-��os�/���0��ʖZJ�
�������Y��s�����;X5��ҳ�m?������/<{tp� U��|-w���q0�Y+`G@�t�门���)Ri����i�o�buʇ앰��ܲ�pm���ri��{�'�h�p`]࡚���p�[
���� �^�Q���+�DR�p ���X:WjϊєĈ��7�Qi�mj]�)JX���E�[��[ �)�n�Sc�W	q�Y�J�>���4����eXo������d�Y�I�\���vX>m �G�P�n58�����N%�Y罒�I��_�O�����+i�(��)��q� "	<�+�x����IPt�a�#�G�A��,�!��>L;}�놢���µ[7ﮑ7�ol{n�����
���7��Q�G��%ky|rR���ds���l$]����+�EV@g��Տ�t:��N5��e�Sc=�mC�֗��Vn �:����w����V�jd�#�Z�P'+**�<������씜����A��a4p�f��a���� 䗣�	����!�BJa�e�9s�	��˥+_f:?7LY��]��!�mӝ,a��m� � ����f�{Y���X��.f�����I�����ݐ+U}Qj_$5Xv���YvCU�ox��:�7�t�_Z�N�yN����nOnT�+.���ѳ[wk{�ue}mm-���]�*C<�o�e��L^����h����Ȧ@�MC餏(���1�+���&ȱ��з��!l�m���1h.���/��s&/��NO�)��g���Eّ���C3�l�O������ƅxC����V�r���L��|$ot �j����墘 3���\M�����B˼g&�QKt�e�2�
4���`+]�?:<�a��ҀCM@�~�dP�k�G�f-��~��k�a��~������LpN�_>KD�s*������?��j��G����f�zf&�d���p��/-��ƿ�_�|ì��#�PK   df�X��p=O  )     jsons/user_defined.json�Y]o�8�+����P�ɾ%�w&�4�lf�b@�T+�#yd�٢��+;���d�n�m_"K:�����s�o��׹������������vQ55�ȳ<���bUt�.�����xpa�{�ח��%�,����
���x���ǣq��BiK�sK�&� �
���Q�	!T�����7�����Y�u��x���oS���m��r��.���±�%S$�,Â E�WX]zO��ټ��U��77q'1aN W������;���TK����|��<�&����i����켪����6�Ww�j1������q�aas�\�;w�ܯ��+���f�Wu��
��>s�˶���v��E�_���E�XQL3
��]S-�k��i���՛��w7�[:�~tG�&��K3[���|1	�>��?ß`ħ|럄O��,/s�ς�<��~�/"�:q�o"�2���<q��oWE�L,�c�f�t�_1�b�@p8B�j�XEy8B�Ę%F��E�����Tc2�"��Of18��"��'��D��a�>����|ɿOf1�L'4�Lq��b�i��݈��,��Ej�p��>���vG�5J�L��Z'r �B}���T��0~��b7/y"��G8,��q.Q����#�0��~�~"f8m��j1BaJ�������kU}�q>�U��;��6s�.�����%���|8�NF���6:#���M���ms�G�}t;���	�z���|��\��6F۲`B i�BF�
i\0Ą�ԃ-*�'Y�{,��D�L��G�%�(�=+y��`)��`Ō���
�!�"f`vI
j�� Z��SD�ᆇ*�q������ၗ4��<{��\�W5<|�/e2����L2���'�i9����9fZ������^`ͲiG���o���G��S΃�n=Gx��e
)�s�UA���G7	1���c���@�%��hn���������ߡ�V�S˛��j�ɑd4���2^�Ӌ��� B����������'Ç'X����,><���aO᯦�ӛ�~�$�>�N�2�� �pj��~_A�^@���j���/�����Cx���.�X{?���`��!n�f 9���`
�~��|0pd}��	�}�XP�|�	�t��B!K�G��Զ�
¼(���x�P��c��?���7'ռ������ڇ�]�m�5Ū�HJ�Qn%C�*�T��<��L�L�����i�)���@�D����v�4����ޏ��
4�}�r��_��UDe����O��<���&(�"���P��/Lr8�q�54����<N�c�@��qeZ�h���بݾ[����Cj����E���,�k��b�{<����m�y>�۰�n^��3[uGt�}˱|�������ȼ͸��m���(�����պ}���[�P4S�Jc��ַ{a��)�U���n��9��i<�]�q�%+��z�X�s���@�a�{*�����.LnG'f����ћ��������V ��%P���,x A$ҮK�*!���H�ڴ��E�F�,�:p�Nq�)0��E�� <����<�+5�[`�}�zV�f�JE�Mpb��9��?��O�'#6�YZrT�050=/+`�7�{��u�df���럫zt�7:�����n>��
�%��\k��z[�R�����Aqi
��0Ҙ/���@�,`�Y�x�RkN3#4U�à� �
T�T�C�d2��0	�Y��v�7��ǿ���1|�>����)}=��%��I_���nOó�"~�<������v���|�,����W��_«߷����$R=��#�H�������f��w{i�}���/�$��'j��������C)=��זGe�mG<�$��Q'��S�#@3I�z�h7���ʻ�����[̌��������:�_�vQ�E�	*qQ gE�;�����HVB���e�ͩ#y�)L.Z�T)»MX!�t)j�f���<�M.�qKx��"���+"��������؟�=xJY&@��h\���ϭ=|֦s6/��i�?����@>��Z����R3�ߠ����:�m�S���B�R-~X�}��_PK
   df�X�xb _  ^�                   cirkitFile.jsonPK
   �b�X�H2�    /             �  images/17766975-adcb-4bce-a273-4a591672b910.pngPK
   6d�X�@M��  2�  /             �'  images/1a44c3f5-ff5c-43a5-9e5f-4b6f5eea1ee8.pngPK
   8f�X\��䓝 Wt /             ��  images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.pngPK
   8f�X���  �  /             �T images/5d57974f-fced-4f10-a93b-7d150e366d9f.pngPK
   tb�X ���s� �� /             q images/5d7124d6-db61-4e16-b8be-eda918c3976e.pngPK
   c�X��{	  -  /             �5 images/62a7f633-b11c-4122-8d1f-7a295c29ca39.pngPK
   �b�Xk���  ��  /             $M images/7b670e17-d5f7-4cb4-b95e-fc2ea835e4f5.pngPK
   tb�X��"�IY eY /             � images/8cf56d13-717b-4162-83ff-adbc9fee247e.pngPK
   8f�Xt`�,s ʉ /             �e images/94a69387-ae01-476e-9716-f0367b107947.pngPK
   c�X<��)�  �  /             �� images/b5e46968-c26e-44e5-9cb6-c624e6f7a7cb.pngPK
   �d�X��'��Z  jk  /              � images/c2c03d23-e153-4716-8f8a-82529ca6767d.pngPK
   6d�X�Rr5�  5 /             GK images/d706f58f-9a00-4cd4-bd85-1d2b1267c556.pngPK
   8f�Xjڎ�]#  X#  /             �� images/f05b9ad5-5094-4ce0-9263-d8ec2a6ced75.pngPK
   �d�X-��R  �W  /             s images/f94c5a85-a3c7-4a52-8d39-8987b87f6a96.pngPK
   df�X��p=O  )               �Z jsons/user_defined.jsonPK      �  =c   